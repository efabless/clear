* NGSPICE file created from top_right_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

.subckt top_right_tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ bottom_width_0_height_0_subtile_0__pin_reg_out_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ bottom_width_0_height_0_subtile_2__pin_inpad_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ ccff_head_0_0 ccff_head_1 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] clk0 gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_dir_0[0]
+ gfpga_pad_io_soc_dir_0[1] gfpga_pad_io_soc_dir_0[2] gfpga_pad_io_soc_dir_0[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_in_0[0]
+ gfpga_pad_io_soc_in_0[1] gfpga_pad_io_soc_in_0[2] gfpga_pad_io_soc_in_0[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] gfpga_pad_io_soc_out_0[0]
+ gfpga_pad_io_soc_out_0[1] gfpga_pad_io_soc_out_0[2] gfpga_pad_io_soc_out_0[3] isol_n
+ left_width_0_height_0_subtile_0__pin_inpad_0_ left_width_0_height_0_subtile_1__pin_inpad_0_
+ left_width_0_height_0_subtile_2__pin_inpad_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ prog_clk prog_reset reset right_width_0_height_0_subtile_0__pin_O_10_ right_width_0_height_0_subtile_0__pin_O_11_
+ right_width_0_height_0_subtile_0__pin_O_12_ right_width_0_height_0_subtile_0__pin_O_13_
+ right_width_0_height_0_subtile_0__pin_O_14_ right_width_0_height_0_subtile_0__pin_O_15_
+ right_width_0_height_0_subtile_0__pin_O_8_ right_width_0_height_0_subtile_0__pin_O_9_
+ sc_in sc_out test_enable top_width_0_height_0_subtile_0__pin_O_0_ top_width_0_height_0_subtile_0__pin_O_1_
+ top_width_0_height_0_subtile_0__pin_O_2_ top_width_0_height_0_subtile_0__pin_O_3_
+ top_width_0_height_0_subtile_0__pin_O_4_ top_width_0_height_0_subtile_0__pin_O_5_
+ top_width_0_height_0_subtile_0__pin_O_6_ top_width_0_height_0_subtile_0__pin_O_7_
+ top_width_0_height_0_subtile_0__pin_cin_0_ top_width_0_height_0_subtile_0__pin_reg_in_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk net758 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__251
+ VGND VGND VPWR VPWR net251 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__251/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2_ net26 cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_44_prog_clk net762 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold340 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold351 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\] VGND VGND VPWR VPWR net711
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold362 cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR net722
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold395 sb_8__8_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold384 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_leaf_53_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold373 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold639_A net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ net429 cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_head VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_55.mux_l1_in_0__A0 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_294_ sb_8__8_.mux_left_track_47.out VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_45.mux_l1_in_1__341 VGND VGND VPWR VPWR net341 sb_8__8_.mux_left_track_45.mux_l1_in_1__341/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_bottom_track_33.mux_l1_in_1_ net309 net6 sb_8__8_.mem_bottom_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net195
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net284 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_2
XFILLER_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net795
+ net179 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ net459 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xhold170 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail VGND VGND VPWR VPWR net530
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold181 cbx_8__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold192 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net552
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ sb_8__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4__A1 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_47.mux_l1_in_0__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3_ sb_8__8_.mux_left_track_29.out net9
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ net444 VGND VGND
+ VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk net661 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net255 net391 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_28_prog_clk net508 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold337_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_13.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__222 VGND VGND VPWR VPWR net222 cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__222/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input55_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
X_329_ net4 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_bottom_track_59.mux_l2_in_0__319 VGND VGND VPWR VPWR net319 sb_8__8_.mux_bottom_track_59.mux_l2_in_0__319/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net458 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_13.out sky130_fd_sc_hd__buf_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_43.mux_l1_in_0_ net162 net62 sb_8__8_.mem_left_track_43.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk net503 net185 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold621_A cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output161_A net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_55.mux_l2_in_0_ net347 sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_55.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_55.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk
+ net863 net169 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_55.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_91_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2_ net14 sb_8__8_.mux_left_track_39.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_3.mux_l3_in_0_ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA__312__A sb_8__8_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout192_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__A0 sb_8__8_.mux_left_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xhold30 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND
+ VPWR VPWR net390 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold41 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X VGND VGND
+ VPWR VPWR net401 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold74 chany_bottom_in[9] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold63 cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold52 cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold85 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold96 cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X VGND VGND VPWR
+ VPWR net456 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk net653 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out
+ net22 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_1_ net6 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_5 net347 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_47.mux_l1_in_1__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__307__A sb_8__8_.mux_left_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_1.mux_l1_in_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net270 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xhold500 sb_8__8_.mem_left_track_57.mem_out\[0\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold511 sb_8__8_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold533 cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\] VGND VGND VPWR VPWR net893
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold522 sb_8__8_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold544 cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR net904
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_fanout205_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold555 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold588 cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR net948
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold577 sb_8__8_.mem_bottom_track_9.mem_out\[1\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold566 cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net926
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold599 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR net959
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net274 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__mux2_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__A1 sb_8__8_.mux_left_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_15.mux_l1_in_1__325 VGND VGND VPWR VPWR net325 sb_8__8_.mux_left_track_15.mux_l1_in_1__325/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4__A0 sb_8__8_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput97 net97 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput86 net86 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_29_prog_clk net623 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_3.mux_l2_in_1_ net333 net165 sb_8__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_29_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ net456 cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2__A0 net33 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold330 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold352 sb_8__8_.mem_bottom_track_31.ccff_tail VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold341 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold374 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold396 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold385 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold363 cbx_8__8_.cbx_1__8_.ccff_head VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk net624
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_22_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out net16
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ sb_8__8_.mux_left_track_49.out VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mux_left_track_55.mux_l1_in_0__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net487 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_33.mux_l1_in_0_ net154 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__320__A sb_8__8_.mux_bottom_track_55.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk net500 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_21.mux_l1_in_0__A0 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_45.mux_l2_in_0_ sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net588
+ net179 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xhold171 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_5_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xhold193 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold182 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net542
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ sb_8__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out net455
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__315__A sb_8__8_.mux_left_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_0_ net428 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net700 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk net745 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_1__A0 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_59.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_13.mux_l1_in_0__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input48_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_328_ net32 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net774
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_23.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3_ net241 sb_8__8_.mux_bottom_track_45.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_45.mux_l1_in_1_ net311 net400 sb_8__8_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__S cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__237 VGND VGND VPWR VPWR net237
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3__237/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A0 sb_8__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__291
+ VGND VGND VPWR VPWR net291 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__291/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output154_A net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_55.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk
+ net803 net169 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_55.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_34_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1_ net427 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ net390 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A0 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout185_A net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.out sky130_fd_sc_hd__clkbuf_2
Xhold31 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 net377 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold64 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold53 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X VGND VGND
+ VPWR VPWR net402 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold75 net62 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold97 chany_bottom_in[19] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold86 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk net464 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_46_prog_clk net532 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_6 net347 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_60_prog_clk
+ net920 net170 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__246 VGND VGND VPWR VPWR net246
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__246/LO sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold501 sb_8__8_.mem_left_track_51.ccff_tail VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold545 cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net905
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold534 cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net894
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__323__A sb_8__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold512 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR net872
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold523 cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR net883
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold556 sb_8__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold567 sb_8__8_.mem_bottom_track_35.mem_out\[0\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold578 sb_8__8_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold589 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR net949
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_11.mux_l2_in_1__A1 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_55.mux_l1_in_0_ net160 net56 sb_8__8_.mem_left_track_55.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net577 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput98 net98 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput87 net87 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_29_prog_clk net576 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2_ sb_8__8_.mux_left_track_27.out net10
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_3.mux_l2_in_0_ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold19_A test_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold320 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2__A1 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net706 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold342 cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\] VGND VGND VPWR VPWR net702
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold331 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold353 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk net501
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold375 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold386 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold364 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold397 cby_8__8_.cby_8__8_.mem_right_ipin_11.ccff_tail VGND VGND VPWR VPWR net757
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_292_ sb_8__8_.mux_left_track_51.out VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3_ net246 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_43_prog_clk net633 net185 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk net591 net196 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk net709 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__A1 sb_8__8_.mux_left_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_21.mux_l1_in_0__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_3.mux_l1_in_1_ net162 net159 sb_8__8_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xhold150 sb_8__8_.mem_bottom_track_1.ccff_tail VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold161 sb_8__8_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold194 cbx_8__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold172 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold183 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ sb_8__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk net686 net203 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net273 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_1__A1 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_327_ net31 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net526
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_23.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2_ net60 sb_8__8_.mux_bottom_track_27.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_45.mux_l1_in_0_ net156 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__326__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk
+ net930 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_57.mux_l2_in_0_ net318 sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_57.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net259 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input60_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net522 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout178_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold32 chany_bottom_in[1] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold21 net75 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold10 net366 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold54 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold65 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold43 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net403 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xhold76 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X VGND VGND
+ VPWR VPWR net436 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold98 net43 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold87 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_31_prog_clk net579 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net696 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_60_prog_clk
+ net958 net170 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_1__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xhold502 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold535 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\] VGND VGND VPWR VPWR net895
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold524 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\] VGND VGND VPWR VPWR net884
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold513 sb_8__8_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold568 cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR net928
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold546 sb_8__8_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold557 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net917
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold579 sb_8__8_.mem_bottom_track_11.mem_out\[1\] VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ net692 net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk net990 net189 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk net862 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput99 net99 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
XFILLER_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput88 net88 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_29_prog_clk net595 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_57.out sky130_fd_sc_hd__clkbuf_2
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_49.mux_l1_in_1__A1 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__S cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net256 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__mux2_8
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout210_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__334__A sb_8__8_.mux_bottom_track_27.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold310 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk net849 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold321 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net681
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold343 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold332 sb_8__8_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold376 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold365 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold354 cby_8__8_.cby_8__8_.mem_right_ipin_2.ccff_tail VGND VGND VPWR VPWR net714
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold387 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_59.mux_l1_in_0__A0 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold398 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ sb_8__8_.mux_left_track_53.out VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_43_prog_clk net466 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_13.mux_l2_in_0_ sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__329__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_19.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_3.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net54 sb_8__8_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold151 cby_8__8_.ccff_tail VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold140 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold162 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold184 sb_8__8_.mem_left_track_9.mem_out\[1\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold173 sb_8__8_.mem_bottom_track_57.mem_out\[0\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold195 sb_8__8_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_5.mux_l2_in_1__314 VGND VGND VPWR VPWR net314 sb_8__8_.mux_bottom_track_5.mux_l2_in_1__314/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ net682 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_343_ sb_8__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_17.mux_l1_in_0__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_13.mux_l1_in_1_ net324 net163 sb_8__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_326_ net30 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1_ net40 cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__342__A sb_8__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_59_prog_clk
+ net963 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input53_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__S cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_309_ sb_8__8_.mux_left_track_17.out VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net474 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__337__A sb_8__8_.mux_bottom_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net882
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold22 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold11 net991 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 net44 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold55 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xhold77 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X VGND VGND
+ VPWR VPWR net437 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold66 chanx_left_in[10] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold99 cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X VGND VGND
+ VPWR VPWR net459 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold88 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_90_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_34_prog_clk net631 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2_ sb_8__8_.mux_bottom_track_15.out
+ net47 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk net938
+ net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_8 chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net81 net71 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ net909 net170 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_1__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3_ net355 sb_8__8_.mux_left_track_55.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_57.mux_l1_in_0_ net388 net154 sb_8__8_.mem_bottom_track_57.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_57.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xhold514 cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR net874
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold536 sb_8__8_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold525 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\] VGND VGND VPWR VPWR net885
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold503 sb_8__8_.mem_bottom_track_55.mem_out\[0\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_0__A0 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold547 sb_8__8_.mem_bottom_track_59.mem_out\[0\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold558 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR net918
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold569 cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR net929
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net802 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout190_A net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net413 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_7.mux_l2_in_1__350 VGND VGND VPWR VPWR net350 sb_8__8_.mux_left_track_7.mux_l2_in_1__350/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput89 net89 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput78 net78 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_29_prog_clk net586 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk net708 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk
+ net885 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_1_0__f_clk0_A clknet_0_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold311 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold300 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold333 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold344 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold322 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net682
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold355 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold377 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold366 cby_8__8_.cby_8__8_.mem_right_ipin_5.ccff_tail VGND VGND VPWR VPWR net726
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold388 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_bottom_track_59.mux_l1_in_0__A1 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold399 sb_8__8_.mem_left_track_15.ccff_tail VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_85_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_left_track_15.mux_l1_in_1__A1 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold248_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_290_ sb_8__8_.mux_left_track_55.out VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2__A0 net400 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4_ sb_8__8_.mux_left_track_43.out
+ net31 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output122_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_41_prog_clk net660 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_25.mux_l1_in_0__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_11.mux_l2_in_1__323 VGND VGND VPWR VPWR net323 sb_8__8_.mux_left_track_11.mux_l2_in_1__323/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk net648 net183 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_67_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__345__A sb_8__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2__A1 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold152 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold130 cby_8__8_.cby_8__8_.mem_right_ipin_3.ccff_tail VGND VGND VPWR VPWR net490
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold141 sb_8__8_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold174 cby_8__8_.cby_8__8_.mem_left_ipin_2.ccff_tail VGND VGND VPWR VPWR net534
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold163 cby_8__8_.cby_8__8_.mem_left_ipin_3.ccff_tail VGND VGND VPWR VPWR net523
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold185 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\] VGND VGND VPWR VPWR net545
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold196 sb_8__8_.mem_bottom_track_25.mem_out\[0\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__282
+ VGND VGND VPWR VPWR net282 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__282/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_18_prog_clk net656 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold365_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ net784 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_342_ sb_8__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_17.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_67_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__287
+ VGND VGND VPWR VPWR net287 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__287/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net291 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_31.mux_l1_in_1__334 VGND VGND VPWR VPWR net334 sb_8__8_.mux_left_track_31.mux_l1_in_1__334/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_13.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net49 sb_8__8_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_325_ sb_8__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold91_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_25.mux_l2_in_0_ net330 sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_25.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk
+ net959 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_18_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input46_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__354 VGND VGND VPWR VPWR net354
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__354/LO sky130_fd_sc_hd__conb_1
XFILLER_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_308_ sb_8__8_.mux_left_track_19.out VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk
+ net895 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__sdfrtp_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net790
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold23 net76 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold12 net993 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold45 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold34 cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X VGND VGND
+ VPWR VPWR net394 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xhold78 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net438 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold67 net4 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold89 chanx_left_in[29] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_34_prog_clk net615 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold612_A cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk net834
+ net188 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_9 chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output152_A net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_left_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net850 net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2_ net25 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net295 net448 net80 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xhold526 sb_8__8_.mem_left_track_11.mem_out\[1\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold504 sb_8__8_.mem_left_track_39.ccff_tail VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold515 sb_8__8_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold537 cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR net897
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold548 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net908
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold559 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR net919
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout183_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_29_prog_clk net674 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput79 net79 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net167 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk net558 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_bottom_track_33.mux_l1_in_0__A0 net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk
+ net955 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__277
+ VGND VGND VPWR VPWR net277 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__277/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_27.mux_l2_in_0__331 VGND VGND VPWR VPWR net331 sb_8__8_.mux_left_track_27.mux_l2_in_0__331/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold301 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold312 cby_8__8_.cby_8__8_.mem_right_ipin_4.ccff_tail VGND VGND VPWR VPWR net672
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold334 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR net694
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold323 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold367 cbx_8__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail VGND VGND VPWR VPWR net727
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold378 cby_8__8_.cby_8__8_.mem_right_ipin_8.ccff_tail VGND VGND VPWR VPWR net738
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold345 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR net705
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold356 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold389 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail net71 VGND
+ VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk
+ net925 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__261
+ VGND VGND VPWR VPWR net261 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__261/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3_ sb_8__8_.mux_left_track_31.out
+ net8 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_40_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_39.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk net486
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_39.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_76_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_41_prog_clk net473 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_15.mux_l2_in_0_ net299 sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_15.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output115_A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_25.mux_l1_in_0__A1 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3_ net228 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net370 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk net816 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold142 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold131 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold153 cbx_8__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail VGND VGND VPWR VPWR net513
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold120 sb_8__8_.mem_bottom_track_15.ccff_tail VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold186 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold164 sb_8__8_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold175 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold197 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_18_prog_clk net625 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk net776 net202 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ net694 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ sb_8__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_25.mux_l2_in_0__304 VGND VGND VPWR VPWR net304 sb_8__8_.mux_bottom_track_25.mux_l2_in_0__304/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l2_in_1__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__220 VGND VGND VPWR VPWR net220 cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__220/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_hold642_A net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_324_ sb_8__8_.mux_bottom_track_47.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_19.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold84_A cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ net640 net186 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net523 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_3_ net237 sb_8__8_.mux_bottom_track_47.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input39_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_307_ sb_8__8_.mux_left_track_21.out VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mux_left_track_31.mux_l1_in_1__A1 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk
+ net919 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3_ net356 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xhold13 net995 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold24 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold46 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold35 cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X VGND VGND
+ VPWR VPWR net395 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xhold68 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR
+ VPWR net428 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold57 chany_bottom_in[13] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold79 cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk net637 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ net768 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk net642
+ net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_25.mux_l1_in_0_ net161 net42 sb_8__8_.mem_left_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net493 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold505 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\] VGND VGND VPWR VPWR net865
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold516 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold527 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net887
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold538 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR net898
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold549 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net909
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_hold47_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__D
+ net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk
+ net891 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_37.mux_l2_in_0_ net337 sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_37.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__273
+ VGND VGND VPWR VPWR net273 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__273/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout176_A net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk net622 net201 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__227 VGND VGND VPWR VPWR net227 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__227/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk net596 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_bottom_track_33.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ net980 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l4_in_0_ net443 cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.ccff_tail VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2__A0 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4_ sb_8__8_.mux_left_track_45.out net30
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4__A0 sb_8__8_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold302 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold313 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold324 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold335 sb_8__8_.mem_bottom_track_51.ccff_tail VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold357 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold368 cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\] VGND VGND VPWR VPWR net728
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold346 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold379 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR net739
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk
+ net962 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net293 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__mux2_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2_ sb_8__8_.mux_left_track_19.out
+ net15 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk net677
+ net203 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_49_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_43_prog_clk net470 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_39.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk net611
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_39.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3_ net218 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net447 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold110 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold121 sb_8__8_.mem_left_track_23.ccff_tail VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold143 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold132 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold176 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold165 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR net525
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold154 sb_8__8_.mem_bottom_track_53.mem_out\[0\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold198 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold187 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail VGND VGND VPWR VPWR net547
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_18_prog_clk net483 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_7.mux_l3_in_0_ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net732 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ net714 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_340_ sb_8__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_0__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ net442 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A gfpga_pad_io_soc_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_27.mux_l1_in_0__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ net411 VGND VGND VPWR
+ VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3_ net223 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ net826 net203 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__233 VGND VGND VPWR VPWR net233
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3__233/LO sky130_fd_sc_hd__conb_1
XFILLER_82_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2__A1 sb_8__8_.mux_left_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net571
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_51.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out net5
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_15.mux_l1_in_0_ net16 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold635_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_323_ sb_8__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_27.mux_l2_in_0_ net305 sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_27.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_57.mux_l2_in_0__318 VGND VGND VPWR VPWR net318 sb_8__8_.mux_bottom_track_57.mux_l2_in_0__318/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ net828 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_1__A0 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_19.mux_l1_in_0__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_7.mux_l2_in_1_ net320 net20 sb_8__8_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__D
+ net683 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ net665 net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__235 VGND VGND VPWR VPWR net235
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__235/LO sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_2_ net441 sb_8__8_.mux_bottom_track_35.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk
+ net710 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk
+ net880 net195 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_306_ sb_8__8_.mux_left_track_23.out VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk
+ net867 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__285
+ VGND VGND VPWR VPWR net285 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__285/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.out sky130_fd_sc_hd__clkbuf_2
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2_ net14 cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold14 net77 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold25 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net396 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 chany_bottom_in[14] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xhold69 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X VGND VGND VPWR
+ VPWR net429 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold58 net37 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk net539 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_3.mux_l2_in_1__A1 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__buf_4_0__A cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_15_prog_clk
+ net854 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net188 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net765 net215 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net65 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xhold517 cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\] VGND VGND VPWR VPWR net877
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold506 cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR net866
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold528 sb_8__8_.mem_bottom_track_1.mem_out\[0\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__244 VGND VGND VPWR VPWR net244
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__244/LO sky130_fd_sc_hd__conb_1
Xhold539 cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net899
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk
+ net964 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout169_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_60_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_13.mux_l1_in_1__324 VGND VGND VPWR VPWR net324 sb_8__8_.mux_left_track_13.mux_l1_in_1__324/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ net726 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_27.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_27.out sky130_fd_sc_hd__clkbuf_2
XFILLER_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3_ sb_8__8_.mux_left_track_33.out net7
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold314 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold303 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold325 sb_8__8_.mem_bottom_track_27.mem_out\[0\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold336 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold369 sb_8__8_.mem_left_track_29.ccff_tail VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold347 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold358 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk
+ net647 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out
+ net21 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_35.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk net846
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_41_prog_clk net720 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_15.mux_l2_in_0__299 VGND VGND VPWR VPWR net299 sb_8__8_.mux_bottom_track_15.mux_l2_in_0__299/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_37.mux_l1_in_0_ net159 net36 sb_8__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__D
+ net725 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold100 cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X VGND VGND
+ VPWR VPWR net460 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk net543 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_49.mux_l2_in_0_ sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_49.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout201_A net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold133 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold122 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold144 sb_8__8_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold111 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold177 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold166 sb_8__8_.mem_bottom_track_21.ccff_tail VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold155 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net276 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xhold199 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold188 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_17_prog_clk net564 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net69 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__A1 sb_8__8_.mux_left_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_27.mux_l1_in_0__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_51.mux_l2_in_0_ net345 sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_51.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk
+ net894 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold22_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2_ net28 sb_8__8_.mux_left_track_31.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ net808 net203 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net79 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net524
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out net11
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_59_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_59_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_322_ sb_8__8_.mux_bottom_track_51.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk
+ net900 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk net544
+ net204 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_49.mux_l1_in_1_ net343 net165 sb_8__8_.mem_left_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_1__A1 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_7.mux_l2_in_0_ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout199_A net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_1_ net36 cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ net918 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk
+ net926 net195 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__218 VGND VGND VPWR VPWR net218 cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__218/LO
+ sky130_fd_sc_hd__conb_1
X_305_ sb_8__8_.mux_left_track_25.out VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XANTENNA__293__A sb_8__8_.mux_left_track_49.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk
+ net738 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net179 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__269
+ VGND VGND VPWR VPWR net269 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__269/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold15 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold37 cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold59 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X VGND VGND
+ VPWR VPWR net419 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold48 net38 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkdlybuf4s50_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk
+ net932 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_27.mux_l1_in_0_ net9 net151 sb_8__8_.mem_bottom_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk net860
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_57.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_7.mux_l1_in_1_ net153 net150 sb_8__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_62_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.out sky130_fd_sc_hd__clkbuf_2
Xhold518 cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\] VGND VGND VPWR VPWR net878
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold507 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR net867
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xhold529 cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net889
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_59.mux_l1_in_1__349 VGND VGND VPWR VPWR net349 sb_8__8_.mux_left_track_59.mux_l1_in_1__349/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ net705 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_27.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_43.mux_l1_in_0__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_55.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_55.out sky130_fd_sc_hd__clkbuf_1
XFILLER_88_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net188 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_1__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output150_A net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk
+ net878 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold304 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold315 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold326 cby_8__8_.cby_8__8_.ccff_tail VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold348 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold359 cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_head VGND VGND VPWR VPWR net719
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold337 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk
+ net832 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_11.mux_l2_in_1__297 VGND VGND VPWR VPWR net297 sb_8__8_.mux_bottom_track_11.mux_l2_in_1__297/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net370 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out
+ net24 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_35.mux_l1_in_0__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net575
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[1] sky130_fd_sc_hd__ebufn_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_41_prog_clk net649 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__292
+ VGND VGND VPWR VPWR net292 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__292/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.out sky130_fd_sc_hd__buf_4
XFILLER_94_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net275 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__mux2_4
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4__A0 sb_8__8_.mux_left_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold101 cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X VGND VGND
+ VPWR VPWR net461 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net482 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold123 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold134 sb_8__8_.mem_left_track_27.ccff_tail VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold112 sb_8__8_.mem_bottom_track_17.ccff_tail VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold145 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold167 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold156 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold189 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold178 sb_8__8_.mem_bottom_track_23.ccff_tail VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_18_prog_clk net463 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.out sky130_fd_sc_hd__clkbuf_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_13_prog_clk net693 net197 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk
+ net954 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1_ net8 cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ sb_8__8_.mux_bottom_track_53.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1__A0 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk
+ net981 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk net943
+ net204 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_49.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net59 sb_8__8_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_25.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_43.mux_l2_in_0__340 VGND VGND VPWR VPWR net340 sb_8__8_.mux_left_track_43.mux_l2_in_0__340/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_14_prog_clk net593 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_51.mux_l1_in_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ net58 sb_8__8_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_35.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold640_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_9.mux_l3_in_0_ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net519
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_25.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk
+ net975 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_15_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_304_ sb_8__8_.mux_left_track_27.out VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2_ sb_8__8_.mux_left_track_19.out net15
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ net425 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_51.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_15_prog_clk
+ net893 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
Xhold16 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold27 chanx_left_in[0] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold38 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold49 cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X VGND VGND
+ VPWR VPWR net409 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ net513 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_24_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_19.out sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mem_left_track_57.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net813
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_57.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_7.mux_l1_in_0_ left_width_0_height_0_subtile_3__pin_inpad_0_
+ left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3_ net242 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net254 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xhold508 cby_8__8_.cby_8__8_.mem_right_ipin_1.ccff_tail VGND VGND VPWR VPWR net868
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold519 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\] VGND VGND VPWR VPWR net879
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk
+ net858 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_43.mux_l1_in_0__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_9.mux_l2_in_1_ net351 net165 sb_8__8_.mem_left_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_1__A1 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net265 net433 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA__299__A sb_8__8_.mux_left_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__A1 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk
+ net948 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold305 sb_8__8_.mem_bottom_track_45.ccff_tail VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold316 cbx_8__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold338 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail VGND
+ VGND VPWR VPWR net698 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold349 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold327 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ net855 net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__A1 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout174_A net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4_ net31 net62 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_41_prog_clk net628 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk net616 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_0__S cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold102 cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold113 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold135 sb_8__8_.mem_bottom_track_19.mem_out\[0\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold124 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold146 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold168 sb_8__8_.mem_left_track_57.ccff_tail VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold157 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold179 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_25_prog_clk net582 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_53.mux_l2_in_0_ net316 sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_53.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net188 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_13_prog_clk net550 net197 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk
+ net941 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_0.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[3] sky130_fd_sc_hd__ebufn_8
XFILLER_55_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_53.out sky130_fd_sc_hd__clkbuf_2
X_320_ sb_8__8_.mux_bottom_track_55.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold516_A cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3_ net247 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input67_A gfpga_pad_io_soc_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ net385 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk
+ net646 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__8_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net529
+ net196 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_14_prog_clk net598 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ net797 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net481
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_25.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__352 VGND VGND VPWR VPWR net352
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__352/LO sky130_fd_sc_hd__conb_1
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk
+ net530 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_303_ sb_8__8_.mux_left_track_29.out VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ net412 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_51.mux_l1_in_0__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold75_A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net730 net210 VGND VGND VPWR VPWR cby_8__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_15_prog_clk
+ net966 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold28 net3 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold17 net379 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold39 chanx_left_in[6] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net195
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2_ net56 cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xhold509 cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR net869
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net505 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l4_in_0_ net395 cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_head VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__S cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_9.mux_l2_in_0_ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold429_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_29.mux_l1_in_1__A1 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk
+ net971 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold306 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold317 sb_8__8_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold328 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold339 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ net712 net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold38_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_A net378 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__ebufn_8
Xsb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3_ sb_8__8_.mux_bottom_track_29.out
+ net39 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk net499 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net715 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__D
+ net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__281
+ VGND VGND VPWR VPWR net281 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__281/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ net394 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__255
+ VGND VGND VPWR VPWR net255 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__255/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_9.mux_l1_in_1_ net162 net159 sb_8__8_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_51.mux_l1_in_1__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold103 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold125 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold114 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold136 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold158 sb_8__8_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold147 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold169 sb_8__8_.mem_left_track_7.ccff_tail VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_25_prog_clk net559 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ net386 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net257 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__mux2_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_14_prog_clk net613 net197 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk
+ net541 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__264
+ VGND VGND VPWR VPWR net264 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__264/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net450
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l2_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2_ net393 net32 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net716 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_19.mux_l2_in_0__301 VGND VGND VPWR VPWR net301 sb_8__8_.mux_bottom_track_19.mux_l2_in_0__301/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_14_prog_clk net585 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_11.mux_l3_in_0_ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_53.mux_l1_in_0_ net25 net152 sb_8__8_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_83_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A0 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net167 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout210 net215 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_6
XFILLER_86_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_302_ sb_8__8_.mux_left_track_31.out VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output166_A net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3__A0 sb_8__8_.mux_left_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__D
+ net667 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_15_prog_clk
+ net897 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold29 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold18 net381 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_2
XANTENNA_fanout197_A net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__231 VGND VGND VPWR VPWR net231 cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__231/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_52_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_11.mux_l2_in_1_ net297 net18 sb_8__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net272 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_47.mux_l1_in_0__A0 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net743 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net446 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__225 VGND VGND VPWR VPWR net225 cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__225/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2__A0 net28 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__267
+ VGND VGND VPWR VPWR net267 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__267/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ net461 VGND VGND
+ VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input42_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk
+ net566 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_25.mux_l2_in_0__330 VGND VGND VPWR VPWR net330 sb_8__8_.mux_left_track_25.mux_l2_in_0__330/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold307 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold318 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold329 cbx_8__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail VGND VGND VPWR VPWR net689
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2__A1 net43 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__259
+ VGND VGND VPWR VPWR net259 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__259/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk net572 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk net886
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_19.mux_l2_in_0_ net327 sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_9.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net51 sb_8__8_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold104 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold126 sb_8__8_.mem_left_track_39.mem_out\[0\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold115 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold137 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold148 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold159 sb_8__8_.mem_left_track_25.mem_out\[0\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mux_left_track_21.mux_l2_in_0_ net328 sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__228 VGND VGND VPWR VPWR net228 cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__228/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_bottom_track_23.mux_l2_in_0__303 VGND VGND VPWR VPWR net303 sb_8__8_.mux_bottom_track_23.mux_l2_in_0__303/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mem_left_track_43.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk net540
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_43.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_14_prog_clk net620 net197 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__ebufn_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__357 VGND VGND VPWR VPWR net357 cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__357/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3__A1 net8 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold98_A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__274
+ VGND VGND VPWR VPWR net274 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__274/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_80_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1_ net34 cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net286 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__mux2_4
XFILLER_89_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold490 cby_8__8_.cby_8__8_.mem_left_ipin_1.ccff_tail VGND VGND VPWR VPWR net850
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net618 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_14_prog_clk net654 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_45.mux_l1_in_1__A1 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout211 net215 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_8
Xfanout200 net202 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ sb_8__8_.mux_left_track_33.out VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input72_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_55.mux_l1_in_0__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3__A1 net11 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output159_A net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_1__A0 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_35.mux_l1_in_1__310 VGND VGND VPWR VPWR net310 sb_8__8_.mux_bottom_track_35.mux_l1_in_1__310/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__271
+ VGND VGND VPWR VPWR net271 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__271/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ net621 net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_51.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_13_prog_clk
+ net752 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold19 test_enable VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2_ sb_8__8_.mux_bottom_track_27.out
+ net40 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__279
+ VGND VGND VPWR VPWR net279 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__279/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_23.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_11.mux_l2_in_0_ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_51_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_55.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_47.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__242 VGND VGND VPWR VPWR net242
+ cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_3__242/LO sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l2_in_1__A1 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold80_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_13.mux_l1_in_0__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3__A0 sb_8__8_.mux_left_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input35_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold308 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold319 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__290
+ VGND VGND VPWR VPWR net290 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__290/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_88_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_11.mux_l1_in_1_ net155 net152 sb_8__8_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk net916
+ net203 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk net756 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_29_prog_clk net664 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output141_A net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold105 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold116 cby_8__8_.cby_8__8_.mem_right_ipin_7.ccff_tail VGND VGND VPWR VPWR net476
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold127 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold138 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold149 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_43.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net807
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_43.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_14_prog_clk net609 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__305__A sb_8__8_.mux_left_track_25.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk net775 net185 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_19.mux_l1_in_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ net46 sb_8__8_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_0__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold480 sb_8__8_.mem_bottom_track_59.ccff_tail VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold491 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3_ net229 sb_8__8_.mux_bottom_track_51.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_21.mux_l1_in_0_ net159 net45 sb_8__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_bottom_track_55.mux_l2_in_0__317 VGND VGND VPWR VPWR net317 sb_8__8_.mux_bottom_track_55.mux_l2_in_0__317/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_14_prog_clk net589 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_33.mux_l2_in_0_ sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_33.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout201 net202 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_8
Xfanout212 net215 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_300_ sb_8__8_.mux_left_track_35.out VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_55.mux_l1_in_0__A1 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input65_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_1__A1 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_40_prog_clk net515 net192 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk net875
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net767 net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput1 net999 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_21.mux_l1_in_0__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4_ net32 net34 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold631_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3_ net358 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ net438 VGND VGND VPWR
+ VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ sky130_fd_sc_hd__clkbuf_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_33.mux_l1_in_1_ net335 net165 sb_8__8_.mem_left_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_34_prog_clk net468 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net290 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3_ net238 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__313__A sb_8__8_.mux_left_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_19_prog_clk net839 net202 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_3.mux_l3_in_0_ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_52_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_13.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_49.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__clkbuf_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net261 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__S cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3_ net357 sb_8__8_.mux_left_track_59.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout215_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 gfpga_pad_io_soc_in_0[3] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail net71 VGND
+ VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_11.mux_l1_in_0_ net157 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4_ sb_8__8_.mux_left_track_41.out net32
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_57.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ net533 net169 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_57.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk net778
+ net203 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk net820 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_13.mux_l2_in_0__298 VGND VGND VPWR VPWR net298 sb_8__8_.mux_bottom_track_13.mux_l2_in_0__298/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_28_prog_clk net945 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output134_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_23.mux_l2_in_0_ net303 sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_23.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_3__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xhold117 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold106 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold128 sb_8__8_.mem_left_track_53.mem_out\[0\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold139 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_3.mux_l2_in_1_ net307 net22 sb_8__8_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold640 ccff_head_1 VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_14_prog_clk net502 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk net829 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l2_in_1__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3_ net219 sb_8__8_.mux_left_track_51.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_23.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_23.out sky130_fd_sc_hd__clkbuf_1
XFILLER_89_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold481 sb_8__8_.mem_left_track_41.mem_out\[0\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold470 sb_8__8_.mem_bottom_track_11.ccff_tail VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__263
+ VGND VGND VPWR VPWR net263 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__263/LO
+ sky130_fd_sc_hd__conb_1
Xhold492 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_2_ net57 cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net504
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_14_prog_clk net678 net197 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__316__A sb_8__8_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__359 VGND VGND VPWR VPWR net359 cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__359/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net268 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__mux2_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3__A1 net37 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xfanout202 net216 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_4
Xfanout213 net215 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_8
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ net892 net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net282 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input58_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_39_prog_clk net517 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3_ net224 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net627
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk net475 net187 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__S cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput2 net1003 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.out sky130_fd_sc_hd__clkbuf_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_21.mux_l1_in_0__A1 net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_3_ sb_8__8_.mux_bottom_track_27.out
+ net40 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_57.mux_l1_in_0__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2_ net26 cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output164_A net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_33.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net38 sb_8__8_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_30_prog_clk net639 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold66_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_19_prog_clk net569 net202 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_45.mux_l2_in_0_ sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout195_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ net556 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_25.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4_ sb_8__8_.mux_left_track_45.out net30
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_left_track_49.mux_l1_in_0__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2_ net388 sb_8__8_.mux_left_track_41.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 isol_n VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_4
Xinput60 chany_bottom_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3_ sb_8__8_.mux_left_track_29.out net9
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_57.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk
+ net825 net169 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_57.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_15.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input40_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_45.mux_l1_in_1_ net341 net163 sb_8__8_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold107 cbx_8__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold129 cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\] VGND VGND VPWR VPWR net489
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold118 sb_8__8_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_3.mux_l2_in_0_ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_59_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__319__A sb_8__8_.mux_bottom_track_57.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_3.mux_l2_in_1__307 VGND VGND VPWR VPWR net307 sb_8__8_.mux_bottom_track_3.mux_l2_in_1__307/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold630 net364 VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold641 net987 VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_17_prog_clk net606 net198 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net761 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.ccff_tail net71 VGND
+ VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_49.mux_l1_in_1__313 VGND VGND VPWR VPWR net313 sb_8__8_.mux_bottom_track_49.mux_l1_in_1__313/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_51.out sky130_fd_sc_hd__clkbuf_2
XFILLER_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2_ net27 sb_8__8_.mux_left_track_39.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_23.mux_l1_in_0_ net11 net157 sb_8__8_.mem_bottom_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk net796 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xhold460 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold471 sb_8__8_.mem_left_track_53.ccff_tail VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold482 sb_8__8_.mem_bottom_track_57.ccff_tail VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold493 sb_8__8_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_3.mux_l1_in_1_ net154 net151 sb_8__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__8_.mux_bottom_track_49.mux_l1_in_1__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk net759
+ net178 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_35.mux_l2_in_0_ sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_35.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_14_prog_clk net497 net197 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__A0 sb_8__8_.mux_left_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net741 net215 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xfanout214 net215 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ net552 net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout203 net205 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__A0 sb_8__8_.mux_left_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold402_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xhold290 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.out sky130_fd_sc_hd__buf_4
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_40_prog_clk net471 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2_ net14 cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk net749 net205 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_289_ sb_8__8_.mux_left_track_57.out VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 net387 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__256
+ VGND VGND VPWR VPWR net256 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__256/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4__A0 sb_8__8_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A0 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__327__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2_ sb_8__8_.mux_bottom_track_15.out
+ net47 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold617_A cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_35.mux_l1_in_1_ net310 net5 sb_8__8_.mem_bottom_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input70_A gfpga_pad_io_soc_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_30_prog_clk net604 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output157_A net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk net913
+ net205 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2__A0 sb_8__8_.mux_left_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_1.mux_l1_in_0__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_23.mux_l1_in_0__A0 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout188_A net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net538 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_25.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_39.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_39.out sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3_ sb_8__8_.mux_left_track_33.out net7
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_2
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_38_prog_clk
+ net581 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1_ net32 cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net279 net424 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput72 prog_reset VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xinput50 chany_bottom_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
Xinput61 chany_bottom_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
XANTENNA__340__A sb_8__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out net16
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_1__A0 net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_15.mux_l1_in_0__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net809 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input33_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_45.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net61 sb_8__8_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold108 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__S cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold119 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A0 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__335__A sb_8__8_.mux_bottom_track_25.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_57.mux_l2_in_0_ net348 sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_57.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__249
+ VGND VGND VPWR VPWR net249 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__249/LO
+ sky130_fd_sc_hd__conb_1
Xhold620 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR net980
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold631 sc_in VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold642 net363 VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_15.out sky130_fd_sc_hd__clkbuf_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_17_prog_clk net597 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net736 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_5.mux_l3_in_0_ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2_ sb_8__8_.mux_left_track_23.out net12
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net271 net406 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout170_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1_ net4 cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net583 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold472 cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail VGND VGND VPWR VPWR net832
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold450 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold461 sb_8__8_.mem_left_track_33.ccff_tail VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold494 cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR net854
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold483 sb_8__8_.mem_bottom_track_5.ccff_tail VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_3.mux_l1_in_0_ net156 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3_ net232 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net506 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold89_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xfanout204 net205 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_6
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk
+ net969 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout215 net216 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_5.mux_l2_in_1_ net344 net166 sb_8__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__260
+ VGND VGND VPWR VPWR net260 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__260/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk net603 net201 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold280 sb_8__8_.mem_bottom_track_47.mem_out\[0\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold291 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_32_prog_clk net718 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net250 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__mux2_8
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_288_ sb_8__8_.mux_left_track_59.out VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_8__8_.mux_left_track_31.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ net711 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput4 net426 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_2__A1 sb_8__8_.mux_bottom_track_27.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__343__A sb_8__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_35.mux_l1_in_0_ net155 left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4_ sb_8__8_.mux_bottom_track_45.out
+ net60 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_0_ net453 cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__294
+ VGND VGND VPWR VPWR net294 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__294/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input63_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_30_prog_clk net650 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk net888
+ net205 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__S cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_47.mux_l2_in_0_ sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_47.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_5.mux_l2_in_1__344 VGND VGND VPWR VPWR net344 sb_8__8_.mux_left_track_5.mux_l2_in_1__344/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_left_track_23.mux_l1_in_0__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__223 VGND VGND VPWR VPWR net223 cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__223/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__338__A sb_8__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput160 net160 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold295_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__A1 sb_8__8_.mux_left_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ net770 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 chany_bottom_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xinput51 chany_bottom_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
Xinput73 net368 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
Xinput62 net434 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net452
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_1__A1 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net570 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3_ net243 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_47.mux_l1_in_1_ net312 net28 sb_8__8_.mem_bottom_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk net911
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net370 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net378 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xhold109 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_57.mux_l2_in_0__348 VGND VGND VPWR VPWR net348 sb_8__8_.mux_left_track_57.mux_l2_in_0__348/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk net901
+ net188 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout213_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold621 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net981
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold610 cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net970
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold632 net371 VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold643 net988 VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ net398 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk net754 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ net423 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__272
+ VGND VGND VPWR VPWR net272 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__272/LO
+ sky130_fd_sc_hd__conb_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk
+ net879 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__346__A sb_8__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1__A0 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk
+ net939 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold451 cbx_8__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail VGND VGND VPWR VPWR net811
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold440 cby_8__8_.cby_8__8_.mem_right_ipin_14.ccff_tail VGND VGND VPWR VPWR net800
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold462 sb_8__8_.mem_left_track_17.ccff_tail VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold484 cby_8__8_.cby_8__8_.mem_right_ipin_0.ccff_tail VGND VGND VPWR VPWR net844
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold473 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\] VGND VGND VPWR VPWR net833
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold495 sb_8__8_.mem_bottom_track_33.mem_out\[0\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold542_A cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2_ net44 cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_1__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_bottom_track_17.mux_l2_in_0__300 VGND VGND VPWR VPWR net300 sb_8__8_.mux_bottom_track_17.mux_l2_in_0__300/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_57.mux_l1_in_0_ net161 net55 sb_8__8_.mem_left_track_57.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__289
+ VGND VGND VPWR VPWR net289 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__289/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ net410 cby_8__8_.cby_8__8_.mem_right_ipin_5.ccff_tail VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ net780 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout205 net216 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net72 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_5.mux_l2_in_0_ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net405 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold270 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold281 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold292 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_32_prog_clk net746 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_31.mux_l1_in_0__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ net949 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net383 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3_ sb_8__8_.mux_bottom_track_33.out
+ net37 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk
+ net728 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_30_prog_clk net675 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input56_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk net511
+ net204 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__240 VGND VGND VPWR VPWR net240
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__240/LO sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_5.mux_l1_in_1_ net163 net160 sb_8__8_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_339_ sb_8__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_23.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net431 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_10 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput161 net161 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput150 net150 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold288_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold455_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold622_A cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output162_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__238 VGND VGND VPWR VPWR net238
+ cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_3__238/LO sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ net912 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1__A0 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_19.mux_l1_in_0__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
Xinput63 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3__A0 sb_8__8_.mux_left_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput41 chany_bottom_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput52 chany_bottom_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
Xinput74 net992 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2_ net58 sb_8__8_.mux_bottom_track_31.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_47.mux_l1_in_0_ net157 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_33_prog_clk net563 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__284
+ VGND VGND VPWR VPWR net284 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__284/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_18_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net821
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_1__A0 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_bottom_track_31.mux_l1_in_1__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_59.mux_l2_in_0_ net319 sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_59.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net172
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk net859
+ net188 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xhold600 cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR net960
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold611 cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR net971
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold633 net74 VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold622 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR net982
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ net398 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net469 net202 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_21.mux_l2_in_0__302 VGND VGND VPWR VPWR net302 sb_8__8_.mux_bottom_track_21.mux_l2_in_0__302/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__247 VGND VGND VPWR VPWR net247
+ cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_3__247/LO sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net785 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold27_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_46_prog_clk
+ net951 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ net873 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_59.mux_l1_in_1__A1 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold463 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_8_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold452 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\] VGND VGND VPWR VPWR net812
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold441 sb_8__8_.mem_bottom_track_9.mem_out\[0\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold430 sb_8__8_.mem_left_track_31.ccff_tail VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold485 cbx_8__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold496 cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\] VGND VGND VPWR VPWR net856
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold474 sb_8__8_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_1__A1 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk
+ net883 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ net462 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_0__A0 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout206 net209 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_8
XFILLER_94_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk
+ net865 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold260 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold271 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold293 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold282 sb_8__8_.mem_bottom_track_3.ccff_tail VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_32_prog_clk net643 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_355_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_59.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ net739 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_83_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net252 net375 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold94_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_left_track_17.mux_l1_in_1__A1 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2__A0 net27 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__253
+ VGND VGND VPWR VPWR net253 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__253/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_15.mux_l2_in_0_ sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_15.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk
+ net904 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_30_prog_clk net666 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input49_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3_ net352 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l3_in_0_ net409 cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[2\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_27.mux_l1_in_0__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ sb_8__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_left_track_5.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net53 sb_8__8_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2__A1 net42 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_11 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput151 net151 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net63 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_87_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ net914 net186 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_7_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk
+ net868 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output155_A net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_19.mux_l1_in_0__A1 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput64 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput42 chany_bottom_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 chany_bottom_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
Xinput75 net380 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XANTENNA_hold57_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__D
+ net669 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__360 VGND VGND VPWR VPWR net360 cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__360/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout186_A net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_15.mux_l1_in_1_ net325 net164 sb_8__8_.mem_left_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out
+ net5 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net370 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net378 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_1_ net408 cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_32_prog_clk net662 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk net843
+ net188 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold612 cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR net972
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold601 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net961
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold634 net372 VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold623 net996 VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_14_prog_clk
+ net681 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk
+ net525 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net915 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_95_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net67 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk
+ net898 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk
+ net773 net186 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_2_ sb_8__8_.mux_bottom_track_19.out
+ net45 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xhold420 cby_8__8_.cby_8__8_.mem_left_ipin_0.ccff_tail VGND VGND VPWR VPWR net780
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold453 sb_8__8_.mem_left_track_55.ccff_tail VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold431 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold442 sb_8__8_.mem_bottom_track_27.ccff_tail VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold475 cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\] VGND VGND VPWR VPWR net835
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold464 cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_head VGND VGND VPWR VPWR net824
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold486 sb_8__8_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_0.out sky130_fd_sc_hd__clkbuf_1
Xhold497 sb_8__8_.mem_left_track_55.mem_out\[0\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net171 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_59.mux_l1_in_0_ net24 net155 sb_8__8_.mem_bottom_track_59.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_59.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_53.mux_l2_in_0__316 VGND VGND VPWR VPWR net316 sb_8__8_.mux_bottom_track_53.mux_l2_in_0__316/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ net929 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk net896
+ net196 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_59_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout207 net209 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_2
XFILLER_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net753 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_59_prog_clk
+ net952 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold250 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold261 sb_8__8_.mem_bottom_track_51.mem_out\[0\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold294 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold272 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold283 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_bottom_track_35.mux_l1_in_0__A0 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_32_prog_clk net629 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_354_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk
+ net672 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_39.mux_l2_in_0__338 VGND VGND VPWR VPWR net338 sb_8__8_.mux_left_track_39.mux_l2_in_0__338/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__D
+ net703 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk net527 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2__A1 sb_8__8_.mux_left_track_39.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net287 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__mux2_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk
+ net972 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk
+ net592 net195 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_30_prog_clk net717 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_27.mux_l1_in_0__A1 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_26_prog_clk net607 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A0 sb_8__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk net488
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_337_ sb_8__8_.mux_bottom_track_21.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_12 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_15.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput152 net152 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk
+ net908 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold343_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ net783 net186 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net374 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input61_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l2_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput54 chany_bottom_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
Xinput43 net457 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput65 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xinput76 net382 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_15_prog_clk
+ net889 net198 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout179_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_15.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net48 sb_8__8_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out
+ net11 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_32_prog_clk net594 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_27.mux_l2_in_0_ net331 sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_27.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk net584 net200 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold602 cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR net962
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold635 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net995
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold624 net998 VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold613 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR net973
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_13_prog_clk
+ net924 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net66 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ net398 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk
+ net957 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_33.mux_l1_in_1__A1 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ net476 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__D
+ net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout211_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk net549 net210 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xhold410 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net770
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold421 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold443 sb_8__8_.mem_bottom_track_53.ccff_tail VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold432 sb_8__8_.mem_left_track_23.mem_out\[0\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold454 sb_8__8_.mem_bottom_track_21.mem_out\[0\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold476 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold465 sb_8__8_.mem_bottom_track_55.ccff_tail VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold487 sb_8__8_.mem_bottom_track_3.mem_out\[1\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold498 cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_tail VGND VGND VPWR VPWR net858
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk net737 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk
+ net560 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2__A0 net26 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_35_prog_clk net516 net203 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk net600
+ net196 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout208 net209 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_4
XANTENNA_hold32_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3_ net234 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_26_prog_clk net485 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk
+ net950 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold262 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail VGND
+ VGND VPWR VPWR net622 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold240 sb_8__8_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold251 sb_8__8_.mem_left_track_37.ccff_tail VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold273 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold284 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__clkbuf_1
Xhold295 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_bottom_track_35.mux_l1_in_0__A1 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_32_prog_clk net602 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_353_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net70 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xsb_8__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net555
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net479 net200 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_17.mux_l2_in_0_ net300 sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_17.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk
+ net835 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3_ net230 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk
+ net719 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ net480 net203 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_26_prog_clk net599 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net861
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4_ net31 net62 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_4__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_336_ sb_8__8_.mux_bottom_track_23.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_13 cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput142 net142 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk
+ net887 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net288 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_7.mux_l1_in_0__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_29.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__289__A sb_8__8_.mux_left_track_57.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__A1 net20 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_319_ sb_8__8_.mux_bottom_track_57.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xinput33 chany_bottom_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 chany_bottom_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput44 net392 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput77 net373 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
Xinput66 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_15_prog_clk
+ net905 net198 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_4_ net31 net62 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__355 VGND VGND VPWR VPWR net355
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__355/LO sky130_fd_sc_hd__conb_1
XFILLER_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out
+ net18 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_32_prog_clk net652 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3_ net359 sb_8__8_.mux_left_track_43.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net557 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output160_A net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_1__A0 net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3_ net239 sb_8__8_.mux_bottom_track_51.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_51.mux_l1_in_0__A0 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
Xhold603 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net963
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold636 ccff_head_0_0 VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold614 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net974
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold625 net1 VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_left_track_59.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk net967
+ net174 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.ccff_head sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk
+ net902 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout191_A net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net772 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold201_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk
+ net965 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3_ net220 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_47.mux_l1_in_1__312 VGND VGND VPWR VPWR net312 sb_8__8_.mux_bottom_track_47.mux_l1_in_1__312/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold400 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold411 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold444 sb_8__8_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold433 sb_8__8_.mem_left_track_27.mem_out\[0\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold422 sb_8__8_.mem_bottom_track_29.ccff_tail VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_left_track_5.mux_l2_in_1__A1 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold455 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_8__8_.mux_left_track_27.mux_l1_in_0_ net162 net41 sb_8__8_.mem_left_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xhold477 sb_8__8_.mem_bottom_track_19.ccff_tail VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold466 sb_8__8_.mem_bottom_track_15.mem_out\[0\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold488 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold499 sb_8__8_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk net536 net205 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk
+ net877 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_70_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net414 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__250
+ VGND VGND VPWR VPWR net250 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__250/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mux_left_track_39.mux_l2_in_0_ net338 sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_39.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk
+ net689 net195 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk net794 net203 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__297__A sb_8__8_.mux_left_track_41.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk net805
+ net203 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net195
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout209 net216 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_11_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2_ net56 cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_41.mux_l2_in_0_ net339 sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_41.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_57_prog_clk
+ net824 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold241 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold252 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold230 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold263 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold296 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold285 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold274 sb_8__8_.mem_left_track_25.ccff_tail VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk net484 net207 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out net5
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_352_ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net518
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__254
+ VGND VGND VPWR VPWR net254 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__254/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_57_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk
+ net960 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_37.mux_l1_in_0__A0 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_2_ net56 cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ net430 VGND VGND VPWR
+ VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ sky130_fd_sc_hd__clkbuf_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_2__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_26_prog_clk net659 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3_ sb_8__8_.mux_bottom_track_29.out
+ net39 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
X_335_ sb_8__8_.mux_bottom_track_25.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_bottom_track_9.mux_l3_in_0_ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net269 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__mux2_4
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__221 VGND VGND VPWR VPWR net221 cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__221/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_hold92_A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput110 net110 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk
+ net935 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_29.mux_l1_in_0__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3_ net225 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input47_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_318_ sb_8__8_.mux_bottom_track_59.out VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_bottom_track_17.mux_l1_in_0_ net15 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput45 chany_bottom_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 chany_bottom_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput67 gfpga_pad_io_soc_in_0[0] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput56 chany_bottom_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk net789 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk net793
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_27.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk
+ net838 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_3_ sb_8__8_.mux_bottom_track_29.out
+ net39 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out
+ net21 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_29.mux_l2_in_0_ sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2_ net31 sb_8__8_.mux_left_track_31.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_32_prog_clk net587 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_41.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_41.out sky130_fd_sc_hd__clkbuf_2
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_9.mux_l2_in_1_ net321 net19 sb_8__8_.mem_bottom_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output153_A net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_1__A1 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2_ net57 net32 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_31.mux_l2_in_0_ sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_31.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net188 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__8_.mux_bottom_track_51.mux_l1_in_0__A1 left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_9.mux_l2_in_1__321 VGND VGND VPWR VPWR net321 sb_8__8_.mux_bottom_track_9.mux_l2_in_1__321/LO
+ sky130_fd_sc_hd__conb_1
Xhold615 cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR net975
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold604 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR net964
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold626 net362 VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_left_track_59.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk net528
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_59.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold637 net983 VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_2_prog_clk
+ net723 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout184_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net848 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk
+ net721 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_88_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 net997 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_29.mux_l1_in_1_ net306 net8 sb_8__8_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold401 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1__S cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.out sky130_fd_sc_hd__clkbuf_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold434 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold445 sb_8__8_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold423 sb_8__8_.mem_bottom_track_47.ccff_tail VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold412 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold478 cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net838
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold467 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold456 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_41_prog_clk net670 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xhold489 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_13_prog_clk
+ net928 net197 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__266
+ VGND VGND VPWR VPWR net266 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__266/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_31.mux_l1_in_1_ net308 net7 sb_8__8_.mem_bottom_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ net927 net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net260 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_29.mux_l1_in_1__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4__A0 sb_8__8_.mux_left_track_39.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_51_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_8__8_.mux_left_track_45.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold220 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold253 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold231 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_1__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold242 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold286 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail VGND VGND VPWR VPWR net646
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold275 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 sb_8__8_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold297 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk net707 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out net11
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_351_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__D
+ net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net277 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_67_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk
+ net551 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_37.mux_l1_in_0__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_39.mux_l1_in_0_ net160 net35 sb_8__8_.mem_left_track_39.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net167 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_hold643_A net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_26_prog_clk net671 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_334_ sb_8__8_.mux_bottom_track_27.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_41.mux_l1_in_0_ net161 net34 sb_8__8_.mem_left_track_41.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_41.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__A0 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold85_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_15 chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__276
+ VGND VGND VPWR VPWR net276 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__276/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput100 net100 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
Xsb_8__8_.mux_left_track_53.mux_l2_in_0_ net346 sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_53.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ net568 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_28_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2_ net26 sb_8__8_.mux_left_track_35.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_1.mux_l3_in_0_ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__236 VGND VGND VPWR VPWR net236
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3__236/LO sky130_fd_sc_hd__conb_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_317_ sb_8__8_.mux_left_track_1.out VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput46 chany_bottom_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput35 chany_bottom_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 net449 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xinput68 gfpga_pad_io_soc_in_0[1] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
Xinput57 chany_bottom_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk net851 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_left_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk net634
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_27.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk
+ net676 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2_ sb_8__8_.mux_bottom_track_17.out
+ net46 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out
+ net24 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1_ net8 cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_32_prog_clk net509 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_51.mux_l1_in_1__315 VGND VGND VPWR VPWR net315 sb_8__8_.mux_bottom_track_51.mux_l1_in_1__315/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold439_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_9.mux_l2_in_0_ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_1_ net34 cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout190 net192 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_4
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_55.mux_l2_in_0__347 VGND VGND VPWR VPWR net347 sb_8__8_.mux_left_track_55.mux_l2_in_0__347/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__D
+ net762 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold616 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net976
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold605 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR net965
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold627 net1000 VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_hold48_A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold638 net361 VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__278
+ VGND VGND VPWR VPWR net278 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__278/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout177_A net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_1.mux_l2_in_1_ net322 net164 sb_8__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__245 VGND VGND VPWR VPWR net245
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3__245/LO sky130_fd_sc_hd__conb_1
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_left_track_53.mux_l1_in_0__A0 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 net985 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_29.mux_l1_in_0_ net152 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail net71 VGND
+ VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold402 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold424 cby_8__8_.cby_8__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net784
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold413 sb_8__8_.mem_bottom_track_11.ccff_head VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold435 sb_8__8_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold468 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net828
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold457 cbx_8__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold446 sb_8__8_.mem_left_track_37.mem_out\[0\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold479 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_41_prog_clk net492 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_9.mux_l1_in_1_ net154 net151 sb_8__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_12_prog_clk
+ net874 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_31.mux_l1_in_0_ net153 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net786 net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net699 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_82_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4__A1 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_45.mux_l1_in_0__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold210 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold243 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail VGND
+ VGND VPWR VPWR net603 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_1__A1 net159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold221 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net581
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold232 sb_8__8_.mem_bottom_track_17.mem_out\[0\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold265 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold254 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold287 cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR net647
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold276 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold298 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_57.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_57.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_57.out sky130_fd_sc_hd__buf_4
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_350_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2__A1 net18 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__A1 sb_8__8_.mux_left_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk
+ net798 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__A0 sb_8__8_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_3_ net233 sb_8__8_.mux_bottom_track_59.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold636_A ccff_head_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_26_prog_clk net641 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_333_ sb_8__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net378 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_3.mux_l2_in_1__333 VGND VGND VPWR VPWR net333 sb_8__8_.mux_left_track_3.mux_l2_in_1__333/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4__A1 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__D
+ net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput101 net101 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.out sky130_fd_sc_hd__clkbuf_2
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_1_ net6 cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net251 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__mux2_8
XFILLER_86_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_316_ sb_8__8_.mux_left_track_3.out VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_bottom_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput69 gfpga_pad_io_soc_in_0[2] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
Xinput47 chany_bottom_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
Xinput58 chany_bottom_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_bottom_track_45.mux_l1_in_1__A1 net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__219 VGND VGND VPWR VPWR net219 cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__219/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_31_prog_clk net531 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_27_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input52_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_1__A0 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout180 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_4
Xfanout191 net192 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_6
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4__A0 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_32_prog_clk net512 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_left_track_11.mux_l3_in_0_ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_53.mux_l1_in_0_ net159 net57 sb_8__8_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold606 cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR net966
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold617 cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR net977
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_27.out sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold639 net984 VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold628 net1002 VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__clkbuf_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ net437 cby_8__8_.cby_8__8_.mem_right_ipin_1.ccff_tail VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__283
+ VGND VGND VPWR VPWR net283 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__283/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_1.mux_l2_in_0_ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2_ sb_8__8_.mux_left_track_23.out net12
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold284_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_left_track_53.mux_l1_in_0__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 net1001 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold425 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold436 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold403 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net763
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold414 sb_8__8_.mem_bottom_track_23.mem_out\[0\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold469 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold447 sb_8__8_.mem_left_track_41.ccff_tail VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold458 sb_8__8_.mem_bottom_track_7.ccff_tail VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_40_prog_clk net612 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_9.mux_l1_in_0_ net156 left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3_ net244 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk
+ net554 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net836 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net278 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_11.mux_l2_in_1_ net323 net166 sb_8__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_1.mux_l1_in_1_ net161 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__293
+ VGND VGND VPWR VPWR net293 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__293/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_60_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_60_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold211 sb_8__8_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold200 cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR net560
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold222 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold233 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_fanout202_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold244 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold266 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold255 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold277 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold299 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold288 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail net71 VGND
+ VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_11.mux_l1_in_0__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net249 net384 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4_ sb_8__8_.mux_bottom_track_45.out
+ net60 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net871
+ net175 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk net733 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_2_ net33 net31 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold629_A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_26_prog_clk net614 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_332_ sb_8__8_.mux_bottom_track_31.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ net421 cby_8__8_.cby_8__8_.mem_right_ipin_6.ccff_tail VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_55.mux_l2_in_0_ net317 sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_55.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput102 net102 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[0] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A0 sb_8__8_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net171 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_315_ sb_8__8_.mux_left_track_5.out VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_56_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput37 net417 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput59 net440 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 chany_bottom_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net258 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold90_A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_49.mux_l1_in_1__343 VGND VGND VPWR VPWR net343 sb_8__8_.mux_left_track_49.mux_l1_in_1__343/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net280 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__mux2_4
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ net514 net169 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_53.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_7_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_55.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input45_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_1__A1 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout170 net171 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_8
Xfanout181 net192 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_8
Xfanout192 net72 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_4
XANTENNA_sb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_31_prog_clk net632 net209 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ net439 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0__A1 net24 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold618 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR net978
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold607 sb_8__8_.mem_left_track_59.mem_out\[0\] VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold629 net2 VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out net19
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold611_A cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output151_A net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 net989 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk net787 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold404 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold415 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold426 sb_8__8_.mem_bottom_track_33.ccff_tail VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold437 cby_8__8_.cby_8__8_.mem_right_ipin_13.ccff_tail VGND VGND VPWR VPWR net797
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold459 sb_8__8_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold448 sb_8__8_.mem_bottom_track_13.ccff_tail VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_41_prog_clk net491 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout182_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.out sky130_fd_sc_hd__buf_4
XANTENNA_sb_8__8_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_2_ net393 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_left_track_11.mux_l2_in_0_ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_49.mux_l1_in_0__A0 net150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l3_in_0_ net436 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_1.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net33 sb_8__8_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__D
+ net648 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk net890
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold201 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold223 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold212 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold234 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold278 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold256 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold245 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold267 sb_8__8_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold289 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk net713 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_37.mux_l2_in_0__337 VGND VGND VPWR VPWR net337 sb_8__8_.mux_left_track_37.mux_l2_in_0__337/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net195
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_1__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk net740
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_3_ sb_8__8_.mux_bottom_track_33.out
+ net418 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_11.mux_l1_in_1_ net163 net160 sb_8__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk net766 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_1_ net435 cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_26_prog_clk net630 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_331_ sb_8__8_.mux_bottom_track_33.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__286
+ VGND VGND VPWR VPWR net286 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__286/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_18 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput103 net103 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[1] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_4__A1 net60 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net383 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ net814 net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_314_ sb_8__8_.mux_left_track_7.out VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 net454 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_52_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput49 chany_bottom_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
Xinput38 net407 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__353 VGND VGND VPWR VPWR net353
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__353/LO sky130_fd_sc_hd__conb_1
XANTENNA__314__A sb_8__8_.mux_left_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_2_ sb_8__8_.mux_bottom_track_23.out
+ net42 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3_ net353 sb_8__8_.mux_left_track_51.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_58_prog_clk
+ net695 net171 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l3_in_0_ net420 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[2\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_55.mux_l1_in_0_ net14 net153 sb_8__8_.mem_bottom_track_55.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_55.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2__A1 sb_8__8_.mux_left_track_39.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout171 net179 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_4
Xfanout182 net185 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_6
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout193 net194 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_31_prog_clk net636 net209 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold608 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR net968
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold619 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR net979
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_left_track_47.mux_l1_in_1__A1 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_1__S cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0_ sb_8__8_.mux_left_track_5.out net22
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__309__A sb_8__8_.mux_left_track_17.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net567 net200 VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_38_prog_clk
+ net619 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold5 net367 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk net750 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__S cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold416 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold405 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold427 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold438 cbx_8__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_40_prog_clk net687 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold449 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4_ sb_8__8_.mux_left_track_39.out
+ net4 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__A0 sb_8__8_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_1_ net419 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[0] sky130_fd_sc_hd__ebufn_8
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_41.mux_l2_in_0__339 VGND VGND VPWR VPWR net339 sb_8__8_.mux_left_track_41.mux_l2_in_0__339/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_15.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_49.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_59.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk
+ net907 net170 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_59.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net478
+ net195 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold202 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold235 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold224 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold213 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold246 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold257 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold268 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold279 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk net701 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_15.mux_l1_in_0__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net267 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_2_ sb_8__8_.mux_bottom_track_21.out
+ net43 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_43_prog_clk net655 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__D cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_1__A0 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__317__A sb_8__8_.mux_left_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3__A0 sb_8__8_.mux_left_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__248
+ VGND VGND VPWR VPWR net248 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__248/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_11.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net50 sb_8__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_26_prog_clk net580 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ sb_8__8_.mux_bottom_track_35.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_23.mux_l2_in_0_ net329 sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_23.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input68_A gfpga_pad_io_soc_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput115 net115 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput104 net104 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[2] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_4__S cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk net819
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ net837 net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_313_ sb_8__8_.mux_left_track_9.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput39 chany_bottom_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_4_prog_clk
+ net542 net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_0__A0 net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2_ net27 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout172 net179 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_6
Xfanout183 net185 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_4
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout194 net216 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_4
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_31_prog_clk net657 net209 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold609 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net969
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net262 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__mux2_4
XFILLER_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_25.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__325__A sb_8__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net294 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_57.mux_l1_in_0__A1 net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk
+ net763 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_13.mux_l1_in_1__A1 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2__A0 net31 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input50_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__226 VGND VGND VPWR VPWR net226 cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__226/LO
+ sky130_fd_sc_hd__conb_1
Xhold6 net369 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ net685 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_27.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_45.mux_l1_in_1__311 VGND VGND VPWR VPWR net311 sb_8__8_.mux_bottom_track_45.mux_l1_in_1__311/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold417 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR net777
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold406 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold428 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_40_prog_clk net668 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold439 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold39_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3_ sb_8__8_.mux_left_track_27.out
+ net10 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_23.mux_l1_in_0__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout168_A net370 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_bottom_track_13.mux_l2_in_0_ net298 sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_13.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_bottom_track_59.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk
+ net842 net169 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_59.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold225 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold214 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold203 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold247 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold236 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold258 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold269 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_15.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_8__8_.cby_8__8_.mux_left_ipin_1.out cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out_0[2] sky130_fd_sc_hd__ebufn_8
XFILLER_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ net403 VGND VGND VPWR
+ VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_1_ sb_8__8_.mux_bottom_track_9.out
+ net50 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_43_prog_clk net663 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__229 VGND VGND VPWR VPWR net229 cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l2_in_3__229/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_59_prog_clk
+ net917 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__333__A sb_8__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk net477 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__232 VGND VGND VPWR VPWR net232
+ cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_3__232/LO sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_29.mux_l1_in_1__306 VGND VGND VPWR VPWR net306 sb_8__8_.mux_bottom_track_29.mux_l1_in_1__306/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1__A1 net19 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3_ net235 net30 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__275
+ VGND VGND VPWR VPWR net275 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__275/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput116 net116 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir_0[3] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_48_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__328__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net822
+ net176 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_312_ sb_8__8_.mux_left_track_11.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net195 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__234 VGND VGND VPWR VPWR net234
+ cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_3__234/LO sky130_fd_sc_hd__conb_1
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xinput29 net399 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk
+ net961 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout198_A net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_3_ net231 sb_8__8_.mux_bottom_track_55.out
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_23.mux_l1_in_0_ net160 net43 sb_8__8_.mem_left_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_3.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout173 net179 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout195 net216 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_31_prog_clk net605 net209 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_35.mux_l2_in_0_ sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_35.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__8_.mux_bottom_track_31.mux_l1_in_0__A0 net153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_19.mux_l2_in_0__327 VGND VGND VPWR VPWR net327 sb_8__8_.mux_left_track_19.mux_l2_in_0__327/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net910
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_7.mux_l2_in_1__320 VGND VGND VPWR VPWR net320 sb_8__8_.mux_bottom_track_7.mux_l2_in_1__320/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_14.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__341__A sb_8__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk net847
+ net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_55_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__243 VGND VGND VPWR VPWR net243
+ cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_3__243/LO sky130_fd_sc_hd__conb_1
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk
+ net978 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 reset VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ net769 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_27.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_4_ net30 net61 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_2__S cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold418 sb_8__8_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold407 sb_8__8_.mem_bottom_track_49.ccff_tail VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold429 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_40_prog_clk net578 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__ebufn_8
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2_ sb_8__8_.mux_left_track_15.out
+ net17 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mux_bottom_track_23.mux_l1_in_0__A1 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net167 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3_ net360 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__336__A sb_8__8_.mux_bottom_track_23.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk
+ net833 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_59.mux_l1_in_0__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_35.mux_l1_in_1_ net336 net166 sb_8__8_.mem_left_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold275_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_60_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_left_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_44_prog_clk net815 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_5.mux_l3_in_0_ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold204 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold226 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold215 sb_8__8_.mem_left_track_1.ccff_tail VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold237 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xhold248 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xhold259 cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net619
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__8_.mux_bottom_track_1.mux_l2_in_1__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_35_prog_clk net744 net203 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3_ net221 sb_8__8_.mux_left_track_45.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net285 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0_ sb_8__8_.mux_bottom_track_3.out
+ net53 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_43_prog_clk net691 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_13.mux_l1_in_0_ net17 left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4_ sb_8__8_.mux_left_track_45.out net30
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_59_prog_clk
+ net953 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_17.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_bottom_track_25.mux_l2_in_0_ net304 sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_25.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk net673 net212 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_5.mux_l2_in_1_ net314 net21 sb_8__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xhold590 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR net950
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk net734 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_2_ net61 sb_8__8_.mux_bottom_track_31.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput106 net106 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.out sky130_fd_sc_hd__clkbuf_2
XFILLER_68_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__344__A sb_8__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_23.mux_l2_in_0__329 VGND VGND VPWR VPWR net329 sb_8__8_.mux_left_track_23.mux_l2_in_0__329/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_86_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net171
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__258
+ VGND VGND VPWR VPWR net258 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__258/LO
+ sky130_fd_sc_hd__conb_1
X_311_ sb_8__8_.mux_left_track_13.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 net451 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ net973 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_77_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net283 net416 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_2_ net55 cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__217 VGND VGND VPWR VPWR net217 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__217/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__A sb_8__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__268
+ VGND VGND VPWR VPWR net268 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__268/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk
+ net812 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xfanout174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_6
XANTENNA_sb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net179 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout196 net216 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_4
Xfanout185 net192 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_31_prog_clk net548 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_25.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_25.out sky130_fd_sc_hd__clkbuf_2
XFILLER_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_53.mux_l2_in_0__346 VGND VGND VPWR VPWR net346 sb_8__8_.mux_left_track_53.mux_l2_in_0__346/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__8_.mux_bottom_track_31.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net729
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold81_A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk net933
+ net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__A0 sb_8__8_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3_ net226 sb_8__8_.mux_left_track_49.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk
+ net986 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_35.mux_l1_in_1__336 VGND VGND VPWR VPWR net336 sb_8__8_.mux_left_track_35.mux_l1_in_1__336/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input36_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 net365 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_3_ sb_8__8_.mux_bottom_track_31.out
+ net38 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold408 cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\] VGND VGND VPWR VPWR net768
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold419 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out
+ net20 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_5.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__A0 sb_8__8_.mux_left_track_41.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_35_prog_clk net771 net205 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2_ net14 cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_19.out sky130_fd_sc_hd__clkbuf_2
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk
+ net947 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_35.mux_l1_in_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ net37 sb_8__8_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_59.mux_l1_in_0__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold602_A cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ net389 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2__A0 sb_8__8_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_47.mux_l2_in_0_ sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_47.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_3.mux_l1_in_0__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_44_prog_clk net725 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net378 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_25.mux_l1_in_0__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold216 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold205 sb_8__8_.mem_left_track_35.ccff_tail VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold249 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold238 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4_ sb_8__8_.mux_left_track_37.out net5
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xhold227 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__270
+ VGND VGND VPWR VPWR net270 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__270/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout173_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net806
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3__S cbx_8__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__347__A sb_8__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_33.mux_l1_in_1__309 VGND VGND VPWR VPWR net309 sb_8__8_.mux_bottom_track_33.mux_l1_in_1__309/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk net852 net203 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.out cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2_ net30 sb_8__8_.mux_left_track_27.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_38_prog_clk net937
+ net188 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_43_prog_clk net788 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3_ sb_8__8_.mux_left_track_33.out net7
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_59_prog_clk
+ net974 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_50_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_1__A0 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_17.mux_l1_in_0__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_47.mux_l1_in_1_ net342 net164 sb_8__8_.mem_left_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_5.mux_l2_in_0_ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold580 cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR net940
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold591 cby_8__8_.cby_8__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR net951
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk net546 net201 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_1_ net38 cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput107 net107 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_310_ sb_8__8_.mux_left_track_15.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_left_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk
+ net534 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__8_.mux_left_track_1.mux_l2_in_1__A1 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input66_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ net944 net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_77_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_8__8_.mux_bottom_track_25.mux_l1_in_0_ net10 net150 sb_8__8_.mem_bottom_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
Xsb_8__8_.mux_bottom_track_5.mux_l1_in_1_ net155 net152 sb_8__8_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__355__A cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net172
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk net876 net204 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk
+ net979 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout197 net202 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout175 net179 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_8
Xfanout186 net188 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_8
XFILLER_47_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_34_prog_clk net651 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk
+ net702 net195 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold74_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk net510
+ net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2_ net28 cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net415 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold9 net73 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkdlybuf4s50_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__265
+ VGND VGND VPWR VPWR net265 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__265/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_59_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_47_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_33.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_29_prog_clk net562 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2_ sb_8__8_.mux_bottom_track_19.out
+ net45 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.out sky130_fd_sc_hd__clkbuf_1
Xhold409 sb_8__8_.mem_bottom_track_25.ccff_tail VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out
+ net23 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_35_prog_clk net573 net205 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ net982 net171 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout216_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold428_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold330_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2__A1 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_44_prog_clk net799 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__A1 sb_8__8_.mux_left_track_57.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_25.mux_l1_in_0__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold206 cbx_8__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold217 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold239 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3_ sb_8__8_.mux_left_track_25.out net11
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xhold228 sb_8__8_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__D
+ net690 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk net934
+ net179 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net565
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0__A0 sb_8__8_.mux_left_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 net376 net168 net994 net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1_ net10 cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk net801
+ net186 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2_ sb_8__8_.mux_left_track_21.out net13
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_43_prog_clk net704 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net179
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_23.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold7_A reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk
+ net844 net169 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mux_bottom_track_5.mux_l1_in_1__A1 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net724 net192 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_47.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net60 sb_8__8_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold581 cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR net941
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold570 cby_8__8_.cby_8__8_.mem_right_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net930
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold592 cby_8__8_.cby_8__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR net952
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ net521 net203 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_1.mux_l2_in_1__322 VGND VGND VPWR VPWR net322 sb_8__8_.mux_left_track_1.mux_l2_in_1__322/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_82_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_59.mux_l2_in_0_ sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.ccff_head
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput119 net119 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput108 net108 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput90 net90 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_7.mux_l3_in_0_ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_left_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2_ sb_8__8_.mux_left_track_15.out net17
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk
+ net489 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_17.out sky130_fd_sc_hd__buf_4
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_45_prog_clk net684 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net731 net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk
+ net884 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net445 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net404 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_left_track_47.mux_l1_in_1__342 VGND VGND VPWR VPWR net342 sb_8__8_.mux_left_track_47.mux_l1_in_1__342/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1__A0 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_56_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_5.mux_l1_in_0_ net157 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3_ net240 sb_8__8_.mux_bottom_track_49.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk
+ net777 net173 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l2_in_2__A0 net44 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_left_track_41.mux_l1_in_0__A0 net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout198 net202 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_4
XFILLER_59_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout176 net178 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_8
Xsb_8__8_.mux_left_track_59.mux_l1_in_1_ net349 net166 sb_8__8_.mem_left_track_59.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xfanout187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_34_prog_clk net601 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold625_A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_1__A0 net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__257
+ VGND VGND VPWR VPWR net257 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__257/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_output165_A net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_7.mux_l2_in_1_ net350 net164 sb_8__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk
+ net942 net195 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold67_A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2__A0 sb_8__8_.mux_left_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__D
+ net561 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout196_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_left_track_33.mux_l1_in_0__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net64 cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_30_prog_clk net638 net214 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.ccff_tail net71 VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4_ net4 net35 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net264 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk
+ net490 net176 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout209_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_49.mux_l2_in_0_ sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_49.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk net760 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold323_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_44_prog_clk net703 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output128_A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_54_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_51.mux_l2_in_0_ sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_51.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold207 cbx_8__8_.cbx_1__8_.ccff_tail VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold229 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2_ sb_8__8_.mux_left_track_13.out net18
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xhold218 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_27.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk net853
+ net174 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__280
+ VGND VGND VPWR VPWR net280 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__280/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.out sky130_fd_sc_hd__clkbuf_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk net818
+ net188 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk
+ net881 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_43_prog_clk net635 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l2_in_1__A0 net36 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold90 net24 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk
+ net545 net186 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_3_ net245 sb_8__8_.mux_bottom_track_53.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_49.mux_l1_in_1_ net313 net27 sb_8__8_.mem_bottom_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net68 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR left_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net188 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk net751 net192 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk
+ net899 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold560 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net920
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold571 cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net931
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold582 cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR net942
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold593 cby_8__8_.cby_8__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net953
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_1.mux_l2_in_1__296 VGND VGND VPWR VPWR net296 sb_8__8_.mux_bottom_track_1.mux_l2_in_1__296/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_bottom_track_51.mux_l1_in_1_ net315 net26 sb_8__8_.mem_bottom_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__8_.mux_left_track_17.mux_l1_in_1__326 VGND VGND VPWR VPWR net326 sb_8__8_.mux_left_track_17.mux_l1_in_1__326/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ net830 net203 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l2_in_1__A0 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_33.mux_l1_in_1__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_0.mux_l1_in_3__A1 net37 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput109 net109 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput91 net91 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput80 net80 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XFILLER_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
XFILLER_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold97_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__D
+ net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1_ sb_8__8_.mux_left_track_9.out net20
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk
+ net940 net196 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk net906
+ net196 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_45_prog_clk net680 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold390 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_92_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net175 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk
+ net956 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ net397 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
X_299_ sb_8__8_.mux_left_track_37.out VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_2_ net58 cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ net742 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_41.mux_l1_in_0__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout199 net202 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_8
Xfanout188 net192 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_4
Xsb_8__8_.mux_left_track_59.mux_l1_in_0_ net162 net44 sb_8__8_.mem_left_track_59.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_59.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xfanout177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_6
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_34_prog_clk net617 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1__f_clk0_A clknet_0_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold618_A cby_8__8_.cby_8__8_.mem_left_ipin_0.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_5.mux_l1_in_1__A1 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input71_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_7.mux_l2_in_0_ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_0__A0 net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk
+ net977 net195 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ net495 net177 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__230 VGND VGND VPWR VPWR net230 cby_8__8_.cby_8__8_.mux_left_ipin_2.mux_l2_in_3__230/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2__A1 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk net827 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk net857
+ net169 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_55.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net195
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__224 VGND VGND VPWR VPWR net224 cbx_8__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__224/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_30_prog_clk net688 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_left_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_3_ sb_8__8_.mux_bottom_track_25.out
+ net41 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net281 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__mux2_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk net781 net210 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_7.mux_l1_in_1_ net161 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk
+ net922 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_29.mux_l1_in_0__A0 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_44_prog_clk net683 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input34_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold208 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail VGND VGND VPWR VPWR net568
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1_ sb_8__8_.mux_left_track_7.out net21
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold219 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_9.mux_l1_in_2__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net840
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_66_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ net422 VGND VGND VPWR
+ VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.ccff_tail net71 VGND
+ VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk
+ net921 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_43_prog_clk net658 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold80 chany_bottom_in[6] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold91 chanx_left_in[24] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk
+ net872 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_2_ net56 sb_8__8_.mux_bottom_track_35.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_49.mux_l1_in_0_ net150 left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout171_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__356 VGND VGND VPWR VPWR net356 cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__356/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk
+ net970 net174 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold572 cbx_8__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR net932
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold561 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net921
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold550 sb_8__8_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold594 cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net954
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold583 sb_8__8_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_bottom_track_51.mux_l1_in_0_ net151 left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xoutput81 net81 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput92 net92 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_11.mux_l2_in_3__A1 net30 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0_ sb_8__8_.mux_left_track_3.out net23
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk
+ net870 net196 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net188 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk net936
+ net196 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_45_prog_clk net507 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold380 sb_8__8_.mem_left_track_43.ccff_tail VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold391 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk net810 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__295__A sb_8__8_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk
+ net968 net172 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND
+ VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_298_ sb_8__8_.mux_left_track_39.out VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_17_prog_clk net698 net201 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfrtp_2
Xsb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk net792
+ net171 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_23.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net248 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout167 net378 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_6
Xfanout178 net179 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_4
Xfanout189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_34_prog_clk net779 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net253 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input64_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_bottom_track_9.mux_l1_in_0__A1 left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk
+ net856 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_14_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk
+ net811 net199 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ net472 net187 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk net764 net204 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1__A0 sb_8__8_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_55.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net831
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_55.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__241 VGND VGND VPWR VPWR net241
+ cby_8__8_.cby_8__8_.mux_right_ipin_3.mux_l2_in_3__241/LO sky130_fd_sc_hd__conb_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk net626 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_2_ sb_8__8_.mux_bottom_track_13.out
+ net48 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_17.mux_l2_in_0_ sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_17.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3_ net354 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l3_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__239 VGND VGND VPWR VPWR net239
+ cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_3__239/LO sky130_fd_sc_hd__conb_1
XFILLER_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk net574 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_left_track_7.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net52 sb_8__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold309_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk
+ net869 net193 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_bottom_track_29.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A net444
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_44_prog_clk net561 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A0 net4 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk
+ net923 net176 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_85_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0_ sb_8__8_.mux_left_track_1.out net24
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xhold209 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_29.mux_l1_in_1__332 VGND VGND VPWR VPWR net332 sb_8__8_.mux_left_track_29.mux_l1_in_1__332/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A0 sb_8__8_.mux_bottom_track_19.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout214_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk
+ net976 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_8__8_.mux_bottom_track_7.mux_l2_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__298__A sb_8__8_.mux_left_track_39.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_17.mux_l1_in_1_ net326 net165 sb_8__8_.mem_left_track_17.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xhold70 cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR
+ VPWR net430 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold81 net59 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold92 net19 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4_ sb_8__8_.mux_left_track_41.out
+ net32 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk
+ net946 net181 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_1_ net36 cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_1 net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk net748 net184 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A0 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk
+ net931 net174 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_33_prog_clk net535 net206 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xhold540 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net900
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold562 cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\] VGND VGND VPWR VPWR net922
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold551 sb_8__8_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold595 cby_8__8_.cby_8__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR net955
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold584 sb_8__8_.mem_bottom_track_45.mem_out\[0\] VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold573 sb_8__8_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_4__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__8_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net179 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xoutput82 net82 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput93 net93 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk
+ net727 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk net755
+ net196 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_44_prog_clk net644 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mux_left_track_35.mux_l1_in_1__A1 net166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold370 cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.ccff_tail
+ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold381 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold392 cbx_8__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk net747 net190 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_2_ sb_8__8_.mux_bottom_track_23.out
+ net42 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net167 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_9.out sky130_fd_sc_hd__buf_4
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ net757 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_297_ sb_8__8_.mux_left_track_41.out VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk net520 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mux_bottom_track_45.mux_l1_in_0__A0 net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk net804
+ net171 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_23.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_6.mux_l1_in_0__A1 net53 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout179 net72 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_4
Xfanout168 net370 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_6
XANTENNA_input1_A net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_8__8_.cby_8__8_.mux_left_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_left_ipin_2.out sky130_fd_sc_hd__clkbuf_2
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2__A0 net14 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input57_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk
+ net866 net179 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_349_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_4.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_30_prog_clk net496 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output163_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_1_ sb_8__8_.mux_bottom_track_7.out
+ net51 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2_ net26 cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout194_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_18_prog_clk net735 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__288
+ VGND VGND VPWR VPWR net288 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__288/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_52_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk net903
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_87_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_43_prog_clk net669 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ net782 net178 VGND VGND VPWR VPWR sb_8__8_.mem_bottom_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net263 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__mux2_4
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3__A1 net10 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_3.mux_l1_in_2__A1 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2__S cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net178 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mux_left_track_9.mux_l1_in_0__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk
+ net547 net200 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1__A1 net21 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_17.mux_l1_in_0_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net47 sb_8__8_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xhold71 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold82 cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X VGND VGND
+ VPWR VPWR net442 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold60 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X VGND VGND
+ VPWR VPWR net420 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold93 cbx_8__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X VGND VGND
+ VPWR VPWR net453 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_63_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_30_prog_clk net679 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3_ sb_8__8_.mux_left_track_29.out
+ net9 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ net800 net180 VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l2_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_2 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold28_A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__8_.mux_left_track_29.mux_l2_in_0_ sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_8__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk net823 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l2_in_3__A1 sb_8__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_1.mux_l1_in_4__A1 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk
+ net467 net177 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk net590 net191 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold530 sb_8__8_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold552 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net912
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold563 sb_8__8_.mem_bottom_track_31.mem_out\[0\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold541 sb_8__8_.mem_bottom_track_7.mem_out\[1\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold585 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold596 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR net956
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold574 sb_8__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__8_.mux_left_track_9.mux_l2_in_1__351 VGND VGND VPWR VPWR net351 sb_8__8_.mux_left_track_9.mux_l2_in_1__351/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_31.mux_l2_in_0_ sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_left_track_31.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput94 net94 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput83 net83 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XFILLER_95_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__8_.mux_bottom_track_53.mux_l1_in_0__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__262
+ VGND VGND VPWR VPWR net262 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__262/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__8_.mux_left_track_21.mux_l2_in_0__328 VGND VGND VPWR VPWR net328 sb_8__8_.mux_left_track_21.mux_l2_in_0__328/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_44_prog_clk net667 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold360 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold371 sb_8__8_.mem_bottom_track_35.ccff_tail VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold393 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1__A0 sb_8__8_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold382 cby_8__8_.cby_8__8_.mem_right_ipin_6.ccff_tail VGND VGND VPWR VPWR net742
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__358 VGND VGND VPWR VPWR net358 cbx_8__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__358/LO
+ sky130_fd_sc_hd__conb_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_1_ sb_8__8_.mux_bottom_track_11.out
+ net49 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_296_ sb_8__8_.mux_left_track_43.out VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_29.mux_l1_in_1_ net332 net163 sb_8__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_46_prog_clk net553 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_45.mux_l1_in_0__A1 left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold95_A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__8_.mux_left_track_7.mux_l2_in_1__A1 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net266 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A0 sb_8__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout169 net171 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_4
Xsb_8__8_.mux_left_track_31.mux_l1_in_1_ net334 net164 sb_8__8_.mem_left_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_3_ net236 sb_8__8_.mux_bottom_track_57.out
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xhold190 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mux_left_track_51.mux_l2_in_0__345 VGND VGND VPWR VPWR net345 sb_8__8_.mux_left_track_51.mux_l2_in_0__345/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk
+ net722 net175 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_0__A0 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_348_ cbx_8__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mux_bottom_track_1.mux_l3_in_0_ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_8__8_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__8_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_33.mux_l1_in_1__335 VGND VGND VPWR VPWR net335 sb_8__8_.mux_left_track_33.mux_l1_in_1__335/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_28_prog_clk net610 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold616_A cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_15.mux_l2_in_2__A1 net32 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output156_A net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_19.mux_l2_in_0_ net301 sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_19.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_2.mux_l1_in_0_ sb_8__8_.mux_bottom_track_1.out
+ net54 cby_8__8_.cby_8__8_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net289 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__D
+ net697 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold58_A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_1_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_39.mux_l1_in_0__A0 net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_21.mux_l2_in_0_ net302 sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_bottom_track_21.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_4_ sb_8__8_.mux_bottom_track_45.out
+ net60 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk net494
+ net177 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk
+ net817 net196 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_43_prog_clk net608 net183 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_1.mux_l2_in_1_ net296 net23 sb_8__8_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l4_in_0_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_8__8_.cby_8__8_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_31.mux_l1_in_1__308 VGND VGND VPWR VPWR net308 sb_8__8_.mux_bottom_track_31.mux_l1_in_1__308/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold147_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_21.out sky130_fd_sc_hd__buf_2
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__252
+ VGND VGND VPWR VPWR net252 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__252/LO
+ sky130_fd_sc_hd__conb_1
Xhold50 cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X VGND VGND
+ VPWR VPWR net410 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold72 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold83 cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X VGND VGND
+ VPWR VPWR net443 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold61 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net421 sky130_fd_sc_hd__clkdlybuf4s25_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net292 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__mux2_4
Xhold94 chanx_left_in[21] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_30_prog_clk net465 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2_ sb_8__8_.mux_left_track_17.out
+ net16 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_left_track_23.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net171 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_3 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3_ net217 sb_8__8_.mux_left_track_47.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A0 sb_8__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_60_prog_clk net841
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_41.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__D
+ net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold520 cbx_8__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net880
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold542 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR net902
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold531 cby_8__8_.cby_8__8_.mem_right_ipin_11.mem_out\[2\] VGND VGND VPWR VPWR net891
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold553 sb_8__8_.mem_bottom_track_1.mem_out\[1\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold564 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net924
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold586 cby_8__8_.cby_8__8_.mem_right_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR net946
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold597 cby_8__8_.cby_8__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR net957
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold575 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR net935
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__295
+ VGND VGND VPWR VPWR net295 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__295/LO
+ sky130_fd_sc_hd__conb_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3__A0 sb_8__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_1.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput84 net84 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xoutput95 net95 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_bottom_track_53.mux_l1_in_0__A1 net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l3_in_1_ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_15.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk net791 net189 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net167 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_50_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3_ net222 sb_8__8_.mux_left_track_53.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_44_prog_clk net697 net182 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold350 cby_8__8_.cby_8__8_.mem_right_ipin_14.mem_out\[2\] VGND VGND VPWR VPWR net710
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold361 cby_8__8_.cby_8__8_.mem_right_ipin_12.ccff_tail VGND VGND VPWR VPWR net721
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold383 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold394 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold372 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_8__8_.cby_8__8_.mux_right_ipin_7.mux_l1_in_0_ sb_8__8_.mux_bottom_track_5.out
+ net52 cby_8__8_.cby_8__8_.mem_right_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_364_ net79 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_295_ sb_8__8_.mux_left_track_45.out VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__8_.mux_left_track_29.mux_l1_in_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net40 sb_8__8_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_8__8_.cby_8__8_.mem_left_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net181
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_8__8_.cby_8__8_.mux_left_ipin_0.mux_l1_in_0__A1 net54 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_31.mux_l1_in_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net39 sb_8__8_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l4_in_0_ net402 cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l2_in_2_ net393 cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xhold180 sb_8__8_.mem_left_track_43.mem_out\[0\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold191 cbx_8__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR net551
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1__A0 net427 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ net845 net194 VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__8_.mux_bottom_track_11.mux_l1_in_0__A1 left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__8_.mux_left_track_43.mux_l2_in_0_ net340 sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__8_.mem_left_track_43.ccff_tail VGND VGND VPWR VPWR sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_27.mux_l2_in_0__305 VGND VGND VPWR VPWR net305 sb_8__8_.mux_bottom_track_27.mux_l2_in_0__305/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_347_ sb_8__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net390 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net177 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net168 grid_clb_8__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net167 VGND
+ VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_sb_8__8_.mux_left_track_47.mux_l1_in_0__A0 bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4_ sb_8__8_.mux_left_track_41.out net32
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_28_prog_clk net645 net213 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold609_A cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l4_in_0_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_0_ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__8_.mux_left_track_39.mux_l1_in_0__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ net401 cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_8__8_.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_A
+ cby_8__8_.cby_8__8_.mux_left_ipin_2.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_3_ sb_8__8_.mux_bottom_track_33.out
+ net37 cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net195
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk net690 net185 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_8__8_.mux_bottom_track_1.mux_l2_in_0_ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_87_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4__A0 sb_8__8_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3_ net227 sb_8__8_.mux_left_track_57.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_8__8_.cby_8__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0__S cbx_8__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__8_.mux_bottom_track_19.mux_l1_in_0_ net13 left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__8_.mem_bottom_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold307_A grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_1_ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_8__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xhold40 net29 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xhold73 grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold62 cby_8__8_.cby_8__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X VGND VGND
+ VPWR VPWR net422 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold51 cby_8__8_.cby_8__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net411 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold84 cby_8__8_.cby_8__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X VGND VGND
+ VPWR VPWR net444 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold95 net16 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_90_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_31_prog_clk net498 net208 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1_ sb_8__8_.mux_left_track_11.out
+ net19 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 net339 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2_ net400 sb_8__8_.mux_left_track_35.out
+ cbx_8__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__8_.mux_bottom_track_21.mux_l1_in_0_ net12 net156 sb_8__8_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_8.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ net396 VGND VGND VPWR
+ VPWR cby_8__8_.cby_8__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ sky130_fd_sc_hd__clkbuf_1
Xsb_8__8_.mem_left_track_41.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net864
+ net170 VGND VGND VPWR VPWR sb_8__8_.mem_left_track_41.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__8_.mux_bottom_track_1.mux_l1_in_1_ net153 net150 sb_8__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout212_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold510 cbx_8__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR net870
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold521 cbx_8__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net881
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold532 cby_8__8_.cby_8__8_.mem_left_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net892
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold554 sb_8__8_.mem_bottom_track_49.mem_out\[0\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold543 sb_8__8_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold565 cbx_8__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\] VGND VGND VPWR VPWR net925
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold576 sb_8__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold587 cby_8__8_.cby_8__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR net947
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold598 cby_8__8_.cby_8__8_.mem_left_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net958
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__8_.mux_bottom_track_33.mux_l2_in_0_ sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X sb_8__8_.mem_bottom_track_33.ccff_tail
+ VGND VGND VPWR VPWR sb_8__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_8__8_.cby_8__8_.mux_right_ipin_10.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__8_.mux_left_track_43.sky130_fd_sc_hd__buf_4_0_ sb_8__8_.mux_left_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__8_.mux_left_track_43.out sky130_fd_sc_hd__clkbuf_2
Xoutput85 net85 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput96 net96 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xgrid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_27_prog_clk net537 net211 VGND VGND VPWR VPWR grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_8__8_.cby_8__8_.mux_right_ipin_12.mux_l3_in_0_ net460 cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ cby_8__8_.cby_8__8_.mem_right_ipin_12.mem_out\[2\] VGND VGND VPWR VPWR cby_8__8_.cby_8__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold33_A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

