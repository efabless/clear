magic
tech sky130A
magscale 1 2
timestamp 1679318172
<< obsli1 >>
rect 1104 2159 49864 54417
<< obsm1 >>
rect 1104 1504 50586 54448
<< metal2 >>
rect 1398 56200 1454 57000
rect 4066 56200 4122 57000
rect 6734 56200 6790 57000
rect 9402 56200 9458 57000
rect 12070 56200 12126 57000
rect 14738 56200 14794 57000
rect 17406 56200 17462 57000
rect 20074 56200 20130 57000
rect 22742 56200 22798 57000
rect 25410 56200 25466 57000
rect 28078 56200 28134 57000
rect 30746 56200 30802 57000
rect 33414 56200 33470 57000
rect 36082 56200 36138 57000
rect 38750 56200 38806 57000
rect 41418 56200 41474 57000
rect 44086 56200 44142 57000
rect 46754 56200 46810 57000
rect 49422 56200 49478 57000
rect 1490 0 1546 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 16946 0 17002 800
rect 17682 0 17738 800
rect 18418 0 18474 800
rect 19154 0 19210 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21362 0 21418 800
rect 22098 0 22154 800
rect 22834 0 22890 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25778 0 25834 800
rect 26514 0 26570 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31666 0 31722 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34610 0 34666 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43442 0 43498 800
rect 44178 0 44234 800
rect 44914 0 44970 800
rect 45650 0 45706 800
rect 46386 0 46442 800
rect 47122 0 47178 800
rect 47858 0 47914 800
rect 48594 0 48650 800
<< obsm2 >>
rect 1510 56144 4010 56273
rect 4178 56144 6678 56273
rect 6846 56144 9346 56273
rect 9514 56144 12014 56273
rect 12182 56144 14682 56273
rect 14850 56144 17350 56273
rect 17518 56144 20018 56273
rect 20186 56144 22686 56273
rect 22854 56144 25354 56273
rect 25522 56144 28022 56273
rect 28190 56144 30690 56273
rect 30858 56144 33358 56273
rect 33526 56144 36026 56273
rect 36194 56144 38694 56273
rect 38862 56144 41362 56273
rect 41530 56144 44030 56273
rect 44198 56144 46698 56273
rect 46866 56144 49366 56273
rect 49534 56144 50580 56273
rect 1400 856 50580 56144
rect 1400 711 1434 856
rect 1602 711 2170 856
rect 2338 711 2906 856
rect 3074 711 3642 856
rect 3810 711 4378 856
rect 4546 711 5114 856
rect 5282 711 5850 856
rect 6018 711 6586 856
rect 6754 711 7322 856
rect 7490 711 8058 856
rect 8226 711 8794 856
rect 8962 711 9530 856
rect 9698 711 10266 856
rect 10434 711 11002 856
rect 11170 711 11738 856
rect 11906 711 12474 856
rect 12642 711 13210 856
rect 13378 711 13946 856
rect 14114 711 14682 856
rect 14850 711 15418 856
rect 15586 711 16154 856
rect 16322 711 16890 856
rect 17058 711 17626 856
rect 17794 711 18362 856
rect 18530 711 19098 856
rect 19266 711 19834 856
rect 20002 711 20570 856
rect 20738 711 21306 856
rect 21474 711 22042 856
rect 22210 711 22778 856
rect 22946 711 23514 856
rect 23682 711 24250 856
rect 24418 711 24986 856
rect 25154 711 25722 856
rect 25890 711 26458 856
rect 26626 711 27194 856
rect 27362 711 27930 856
rect 28098 711 28666 856
rect 28834 711 29402 856
rect 29570 711 30138 856
rect 30306 711 30874 856
rect 31042 711 31610 856
rect 31778 711 32346 856
rect 32514 711 33082 856
rect 33250 711 33818 856
rect 33986 711 34554 856
rect 34722 711 35290 856
rect 35458 711 36026 856
rect 36194 711 36762 856
rect 36930 711 37498 856
rect 37666 711 38234 856
rect 38402 711 38970 856
rect 39138 711 39706 856
rect 39874 711 40442 856
rect 40610 711 41178 856
rect 41346 711 41914 856
rect 42082 711 42650 856
rect 42818 711 43386 856
rect 43554 711 44122 856
rect 44290 711 44858 856
rect 45026 711 45594 856
rect 45762 711 46330 856
rect 46498 711 47066 856
rect 47234 711 47802 856
rect 47970 711 48538 856
rect 48706 711 50580 856
<< metal3 >>
rect 50200 56176 51000 56296
rect 50200 55360 51000 55480
rect 50200 54544 51000 54664
rect 50200 53728 51000 53848
rect 50200 52912 51000 53032
rect 50200 52096 51000 52216
rect 50200 51280 51000 51400
rect 50200 50464 51000 50584
rect 50200 49648 51000 49768
rect 50200 48832 51000 48952
rect 50200 48016 51000 48136
rect 50200 47200 51000 47320
rect 50200 46384 51000 46504
rect 50200 45568 51000 45688
rect 50200 44752 51000 44872
rect 50200 43936 51000 44056
rect 50200 43120 51000 43240
rect 50200 42304 51000 42424
rect 50200 41488 51000 41608
rect 50200 40672 51000 40792
rect 50200 39856 51000 39976
rect 50200 39040 51000 39160
rect 50200 38224 51000 38344
rect 50200 37408 51000 37528
rect 50200 36592 51000 36712
rect 50200 35776 51000 35896
rect 50200 34960 51000 35080
rect 50200 34144 51000 34264
rect 50200 33328 51000 33448
rect 50200 32512 51000 32632
rect 50200 31696 51000 31816
rect 50200 30880 51000 31000
rect 50200 30064 51000 30184
rect 50200 29248 51000 29368
rect 50200 28432 51000 28552
rect 50200 27616 51000 27736
rect 50200 26800 51000 26920
rect 50200 25984 51000 26104
rect 50200 25168 51000 25288
rect 50200 24352 51000 24472
rect 50200 23536 51000 23656
rect 50200 22720 51000 22840
rect 50200 21904 51000 22024
rect 50200 21088 51000 21208
rect 50200 20272 51000 20392
rect 50200 19456 51000 19576
rect 50200 18640 51000 18760
rect 50200 17824 51000 17944
rect 50200 17008 51000 17128
rect 50200 16192 51000 16312
rect 50200 15376 51000 15496
rect 50200 14560 51000 14680
rect 50200 13744 51000 13864
rect 50200 12928 51000 13048
rect 50200 12112 51000 12232
rect 50200 11296 51000 11416
rect 50200 10480 51000 10600
rect 50200 9664 51000 9784
rect 0 8712 800 8832
rect 50200 8848 51000 8968
rect 50200 8032 51000 8152
rect 50200 7216 51000 7336
rect 0 6400 800 6520
rect 50200 6400 51000 6520
rect 50200 5584 51000 5704
rect 50200 4768 51000 4888
rect 0 4088 800 4208
rect 50200 3952 51000 4072
rect 50200 3136 51000 3256
rect 50200 2320 51000 2440
rect 0 1776 800 1896
rect 50200 1504 51000 1624
rect 50200 688 51000 808
<< obsm3 >>
rect 800 56096 50120 56269
rect 800 55560 50495 56096
rect 800 55280 50120 55560
rect 800 54744 50495 55280
rect 800 54464 50120 54744
rect 800 53928 50495 54464
rect 800 53648 50120 53928
rect 800 53112 50495 53648
rect 800 52832 50120 53112
rect 800 52296 50495 52832
rect 800 52016 50120 52296
rect 800 51480 50495 52016
rect 800 51200 50120 51480
rect 800 50664 50495 51200
rect 800 50384 50120 50664
rect 800 49848 50495 50384
rect 800 49568 50120 49848
rect 800 49032 50495 49568
rect 800 48752 50120 49032
rect 800 48216 50495 48752
rect 800 47936 50120 48216
rect 800 47400 50495 47936
rect 800 47120 50120 47400
rect 800 46584 50495 47120
rect 800 46304 50120 46584
rect 800 45768 50495 46304
rect 800 45488 50120 45768
rect 800 44952 50495 45488
rect 800 44672 50120 44952
rect 800 44136 50495 44672
rect 800 43856 50120 44136
rect 800 43320 50495 43856
rect 800 43040 50120 43320
rect 800 42504 50495 43040
rect 800 42224 50120 42504
rect 800 41688 50495 42224
rect 800 41408 50120 41688
rect 800 40872 50495 41408
rect 800 40592 50120 40872
rect 800 40056 50495 40592
rect 800 39776 50120 40056
rect 800 39240 50495 39776
rect 800 38960 50120 39240
rect 800 38424 50495 38960
rect 800 38144 50120 38424
rect 800 37608 50495 38144
rect 800 37328 50120 37608
rect 800 36792 50495 37328
rect 800 36512 50120 36792
rect 800 35976 50495 36512
rect 800 35696 50120 35976
rect 800 35160 50495 35696
rect 800 34880 50120 35160
rect 800 34344 50495 34880
rect 800 34064 50120 34344
rect 800 33528 50495 34064
rect 800 33248 50120 33528
rect 800 32712 50495 33248
rect 800 32432 50120 32712
rect 800 31896 50495 32432
rect 800 31616 50120 31896
rect 800 31080 50495 31616
rect 800 30800 50120 31080
rect 800 30264 50495 30800
rect 800 29984 50120 30264
rect 800 29448 50495 29984
rect 800 29168 50120 29448
rect 800 28632 50495 29168
rect 800 28352 50120 28632
rect 800 27816 50495 28352
rect 800 27536 50120 27816
rect 800 27000 50495 27536
rect 800 26720 50120 27000
rect 800 26184 50495 26720
rect 800 25904 50120 26184
rect 800 25368 50495 25904
rect 800 25088 50120 25368
rect 800 24552 50495 25088
rect 800 24272 50120 24552
rect 800 23736 50495 24272
rect 800 23456 50120 23736
rect 800 22920 50495 23456
rect 800 22640 50120 22920
rect 800 22104 50495 22640
rect 800 21824 50120 22104
rect 800 21288 50495 21824
rect 800 21008 50120 21288
rect 800 20472 50495 21008
rect 800 20192 50120 20472
rect 800 19656 50495 20192
rect 800 19376 50120 19656
rect 800 18840 50495 19376
rect 800 18560 50120 18840
rect 800 18024 50495 18560
rect 800 17744 50120 18024
rect 800 17208 50495 17744
rect 800 16928 50120 17208
rect 800 16392 50495 16928
rect 800 16112 50120 16392
rect 800 15576 50495 16112
rect 800 15296 50120 15576
rect 800 14760 50495 15296
rect 800 14480 50120 14760
rect 800 13944 50495 14480
rect 800 13664 50120 13944
rect 800 13128 50495 13664
rect 800 12848 50120 13128
rect 800 12312 50495 12848
rect 800 12032 50120 12312
rect 800 11496 50495 12032
rect 800 11216 50120 11496
rect 800 10680 50495 11216
rect 800 10400 50120 10680
rect 800 9864 50495 10400
rect 800 9584 50120 9864
rect 800 9048 50495 9584
rect 800 8912 50120 9048
rect 880 8768 50120 8912
rect 880 8632 50495 8768
rect 800 8232 50495 8632
rect 800 7952 50120 8232
rect 800 7416 50495 7952
rect 800 7136 50120 7416
rect 800 6600 50495 7136
rect 880 6320 50120 6600
rect 800 5784 50495 6320
rect 800 5504 50120 5784
rect 800 4968 50495 5504
rect 800 4688 50120 4968
rect 800 4288 50495 4688
rect 880 4152 50495 4288
rect 880 4008 50120 4152
rect 800 3872 50120 4008
rect 800 3336 50495 3872
rect 800 3056 50120 3336
rect 800 2520 50495 3056
rect 800 2240 50120 2520
rect 800 1976 50495 2240
rect 880 1704 50495 1976
rect 880 1696 50120 1704
rect 800 1424 50120 1696
rect 800 888 50495 1424
rect 800 715 50120 888
<< metal4 >>
rect 2944 2128 3264 54448
rect 7944 2128 8264 54448
rect 12944 2128 13264 54448
rect 17944 2128 18264 54448
rect 22944 2128 23264 54448
rect 27944 2128 28264 54448
rect 32944 2128 33264 54448
rect 37944 2128 38264 54448
rect 42944 2128 43264 54448
rect 47944 2128 48264 54448
<< obsm4 >>
rect 26006 2347 27864 33693
rect 28344 2347 32864 33693
rect 33344 2347 37661 33693
<< labels >>
rlabel metal4 s 7944 2128 8264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27944 2128 28264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37944 2128 38264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47944 2128 48264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 32944 2128 33264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 42944 2128 43264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 49422 56200 49478 57000 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 ccff_head_0
port 4 nsew signal input
rlabel metal3 s 50200 688 51000 808 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 1398 56200 1454 57000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 50200 25984 51000 26104 6 chanx_right_in[0]
port 7 nsew signal input
rlabel metal3 s 50200 34144 51000 34264 6 chanx_right_in[10]
port 8 nsew signal input
rlabel metal3 s 50200 34960 51000 35080 6 chanx_right_in[11]
port 9 nsew signal input
rlabel metal3 s 50200 35776 51000 35896 6 chanx_right_in[12]
port 10 nsew signal input
rlabel metal3 s 50200 36592 51000 36712 6 chanx_right_in[13]
port 11 nsew signal input
rlabel metal3 s 50200 37408 51000 37528 6 chanx_right_in[14]
port 12 nsew signal input
rlabel metal3 s 50200 38224 51000 38344 6 chanx_right_in[15]
port 13 nsew signal input
rlabel metal3 s 50200 39040 51000 39160 6 chanx_right_in[16]
port 14 nsew signal input
rlabel metal3 s 50200 39856 51000 39976 6 chanx_right_in[17]
port 15 nsew signal input
rlabel metal3 s 50200 40672 51000 40792 6 chanx_right_in[18]
port 16 nsew signal input
rlabel metal3 s 50200 41488 51000 41608 6 chanx_right_in[19]
port 17 nsew signal input
rlabel metal3 s 50200 26800 51000 26920 6 chanx_right_in[1]
port 18 nsew signal input
rlabel metal3 s 50200 42304 51000 42424 6 chanx_right_in[20]
port 19 nsew signal input
rlabel metal3 s 50200 43120 51000 43240 6 chanx_right_in[21]
port 20 nsew signal input
rlabel metal3 s 50200 43936 51000 44056 6 chanx_right_in[22]
port 21 nsew signal input
rlabel metal3 s 50200 44752 51000 44872 6 chanx_right_in[23]
port 22 nsew signal input
rlabel metal3 s 50200 45568 51000 45688 6 chanx_right_in[24]
port 23 nsew signal input
rlabel metal3 s 50200 46384 51000 46504 6 chanx_right_in[25]
port 24 nsew signal input
rlabel metal3 s 50200 47200 51000 47320 6 chanx_right_in[26]
port 25 nsew signal input
rlabel metal3 s 50200 48016 51000 48136 6 chanx_right_in[27]
port 26 nsew signal input
rlabel metal3 s 50200 48832 51000 48952 6 chanx_right_in[28]
port 27 nsew signal input
rlabel metal3 s 50200 49648 51000 49768 6 chanx_right_in[29]
port 28 nsew signal input
rlabel metal3 s 50200 27616 51000 27736 6 chanx_right_in[2]
port 29 nsew signal input
rlabel metal3 s 50200 28432 51000 28552 6 chanx_right_in[3]
port 30 nsew signal input
rlabel metal3 s 50200 29248 51000 29368 6 chanx_right_in[4]
port 31 nsew signal input
rlabel metal3 s 50200 30064 51000 30184 6 chanx_right_in[5]
port 32 nsew signal input
rlabel metal3 s 50200 30880 51000 31000 6 chanx_right_in[6]
port 33 nsew signal input
rlabel metal3 s 50200 31696 51000 31816 6 chanx_right_in[7]
port 34 nsew signal input
rlabel metal3 s 50200 32512 51000 32632 6 chanx_right_in[8]
port 35 nsew signal input
rlabel metal3 s 50200 33328 51000 33448 6 chanx_right_in[9]
port 36 nsew signal input
rlabel metal3 s 50200 1504 51000 1624 6 chanx_right_out[0]
port 37 nsew signal output
rlabel metal3 s 50200 9664 51000 9784 6 chanx_right_out[10]
port 38 nsew signal output
rlabel metal3 s 50200 10480 51000 10600 6 chanx_right_out[11]
port 39 nsew signal output
rlabel metal3 s 50200 11296 51000 11416 6 chanx_right_out[12]
port 40 nsew signal output
rlabel metal3 s 50200 12112 51000 12232 6 chanx_right_out[13]
port 41 nsew signal output
rlabel metal3 s 50200 12928 51000 13048 6 chanx_right_out[14]
port 42 nsew signal output
rlabel metal3 s 50200 13744 51000 13864 6 chanx_right_out[15]
port 43 nsew signal output
rlabel metal3 s 50200 14560 51000 14680 6 chanx_right_out[16]
port 44 nsew signal output
rlabel metal3 s 50200 15376 51000 15496 6 chanx_right_out[17]
port 45 nsew signal output
rlabel metal3 s 50200 16192 51000 16312 6 chanx_right_out[18]
port 46 nsew signal output
rlabel metal3 s 50200 17008 51000 17128 6 chanx_right_out[19]
port 47 nsew signal output
rlabel metal3 s 50200 2320 51000 2440 6 chanx_right_out[1]
port 48 nsew signal output
rlabel metal3 s 50200 17824 51000 17944 6 chanx_right_out[20]
port 49 nsew signal output
rlabel metal3 s 50200 18640 51000 18760 6 chanx_right_out[21]
port 50 nsew signal output
rlabel metal3 s 50200 19456 51000 19576 6 chanx_right_out[22]
port 51 nsew signal output
rlabel metal3 s 50200 20272 51000 20392 6 chanx_right_out[23]
port 52 nsew signal output
rlabel metal3 s 50200 21088 51000 21208 6 chanx_right_out[24]
port 53 nsew signal output
rlabel metal3 s 50200 21904 51000 22024 6 chanx_right_out[25]
port 54 nsew signal output
rlabel metal3 s 50200 22720 51000 22840 6 chanx_right_out[26]
port 55 nsew signal output
rlabel metal3 s 50200 23536 51000 23656 6 chanx_right_out[27]
port 56 nsew signal output
rlabel metal3 s 50200 24352 51000 24472 6 chanx_right_out[28]
port 57 nsew signal output
rlabel metal3 s 50200 25168 51000 25288 6 chanx_right_out[29]
port 58 nsew signal output
rlabel metal3 s 50200 3136 51000 3256 6 chanx_right_out[2]
port 59 nsew signal output
rlabel metal3 s 50200 3952 51000 4072 6 chanx_right_out[3]
port 60 nsew signal output
rlabel metal3 s 50200 4768 51000 4888 6 chanx_right_out[4]
port 61 nsew signal output
rlabel metal3 s 50200 5584 51000 5704 6 chanx_right_out[5]
port 62 nsew signal output
rlabel metal3 s 50200 6400 51000 6520 6 chanx_right_out[6]
port 63 nsew signal output
rlabel metal3 s 50200 7216 51000 7336 6 chanx_right_out[7]
port 64 nsew signal output
rlabel metal3 s 50200 8032 51000 8152 6 chanx_right_out[8]
port 65 nsew signal output
rlabel metal3 s 50200 8848 51000 8968 6 chanx_right_out[9]
port 66 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_in_0[0]
port 67 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in_0[10]
port 68 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in_0[11]
port 69 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in_0[12]
port 70 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in_0[13]
port 71 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_in_0[14]
port 72 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_in_0[15]
port 73 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_in_0[16]
port 74 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_in_0[17]
port 75 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_in_0[18]
port 76 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 chany_bottom_in_0[19]
port 77 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 chany_bottom_in_0[1]
port 78 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_in_0[20]
port 79 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_in_0[21]
port 80 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_in_0[22]
port 81 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_in_0[23]
port 82 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_in_0[24]
port 83 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_in_0[25]
port 84 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_in_0[26]
port 85 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_in_0[27]
port 86 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 chany_bottom_in_0[28]
port 87 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 chany_bottom_in_0[29]
port 88 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in_0[2]
port 89 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_in_0[3]
port 90 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in_0[4]
port 91 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in_0[5]
port 92 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in_0[6]
port 93 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in_0[7]
port 94 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in_0[8]
port 95 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in_0[9]
port 96 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 chany_bottom_out_0[0]
port 97 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 chany_bottom_out_0[10]
port 98 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 chany_bottom_out_0[11]
port 99 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 chany_bottom_out_0[12]
port 100 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 chany_bottom_out_0[13]
port 101 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 chany_bottom_out_0[14]
port 102 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 chany_bottom_out_0[15]
port 103 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 chany_bottom_out_0[16]
port 104 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 chany_bottom_out_0[17]
port 105 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 chany_bottom_out_0[18]
port 106 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 chany_bottom_out_0[19]
port 107 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 chany_bottom_out_0[1]
port 108 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 chany_bottom_out_0[20]
port 109 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 chany_bottom_out_0[21]
port 110 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 chany_bottom_out_0[22]
port 111 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 chany_bottom_out_0[23]
port 112 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 chany_bottom_out_0[24]
port 113 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 chany_bottom_out_0[25]
port 114 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 chany_bottom_out_0[26]
port 115 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 chany_bottom_out_0[27]
port 116 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 chany_bottom_out_0[28]
port 117 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 chany_bottom_out_0[29]
port 118 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 chany_bottom_out_0[2]
port 119 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 chany_bottom_out_0[3]
port 120 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 chany_bottom_out_0[4]
port 121 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 chany_bottom_out_0[5]
port 122 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 chany_bottom_out_0[6]
port 123 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 chany_bottom_out_0[7]
port 124 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 chany_bottom_out_0[8]
port 125 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 chany_bottom_out_0[9]
port 126 nsew signal output
rlabel metal2 s 4066 56200 4122 57000 6 gfpga_pad_io_soc_dir[0]
port 127 nsew signal output
rlabel metal2 s 6734 56200 6790 57000 6 gfpga_pad_io_soc_dir[1]
port 128 nsew signal output
rlabel metal2 s 9402 56200 9458 57000 6 gfpga_pad_io_soc_dir[2]
port 129 nsew signal output
rlabel metal2 s 12070 56200 12126 57000 6 gfpga_pad_io_soc_dir[3]
port 130 nsew signal output
rlabel metal2 s 25410 56200 25466 57000 6 gfpga_pad_io_soc_in[0]
port 131 nsew signal input
rlabel metal2 s 28078 56200 28134 57000 6 gfpga_pad_io_soc_in[1]
port 132 nsew signal input
rlabel metal2 s 30746 56200 30802 57000 6 gfpga_pad_io_soc_in[2]
port 133 nsew signal input
rlabel metal2 s 33414 56200 33470 57000 6 gfpga_pad_io_soc_in[3]
port 134 nsew signal input
rlabel metal2 s 14738 56200 14794 57000 6 gfpga_pad_io_soc_out[0]
port 135 nsew signal output
rlabel metal2 s 17406 56200 17462 57000 6 gfpga_pad_io_soc_out[1]
port 136 nsew signal output
rlabel metal2 s 20074 56200 20130 57000 6 gfpga_pad_io_soc_out[2]
port 137 nsew signal output
rlabel metal2 s 22742 56200 22798 57000 6 gfpga_pad_io_soc_out[3]
port 138 nsew signal output
rlabel metal2 s 36082 56200 36138 57000 6 isol_n
port 139 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 prog_clk
port 140 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 prog_reset_bottom_in
port 141 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 reset_bottom_in
port 142 nsew signal input
rlabel metal3 s 50200 50464 51000 50584 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 143 nsew signal input
rlabel metal3 s 50200 51280 51000 51400 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 144 nsew signal input
rlabel metal3 s 50200 52096 51000 52216 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 145 nsew signal input
rlabel metal3 s 50200 52912 51000 53032 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 146 nsew signal input
rlabel metal3 s 50200 53728 51000 53848 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 147 nsew signal input
rlabel metal3 s 50200 54544 51000 54664 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 148 nsew signal input
rlabel metal3 s 50200 55360 51000 55480 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 149 nsew signal input
rlabel metal3 s 50200 56176 51000 56296 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 150 nsew signal input
rlabel metal2 s 38750 56200 38806 57000 6 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
rlabel metal2 s 41418 56200 41474 57000 6 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
rlabel metal2 s 44086 56200 44142 57000 6 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
rlabel metal2 s 46754 56200 46810 57000 6 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 right_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 right_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 right_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 right_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 test_enable_bottom_in
port 159 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51000 57000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2493530
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/top_left_tile/runs/23_03_20_06_14/results/signoff/top_left_tile.magic.gds
string GDS_START 170388
<< end >>

