VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2475.000 BY 2715.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -12.760 -3.720 -7.960 2718.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 -3.720 2487.560 1.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2713.480 2487.560 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2482.760 -3.720 2487.560 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.920 -3.720 13.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 -3.720 70.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 174.765 70.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 477.540 70.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 792.540 70.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 1107.540 70.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 1422.540 70.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 1737.540 70.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 2052.540 70.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 2367.540 70.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.920 2682.540 70.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 -3.720 127.120 45.715 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 174.765 127.120 200.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 475.085 127.120 515.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 790.085 127.120 830.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 1105.085 127.120 1145.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 1420.085 127.120 1460.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 1735.085 127.120 1775.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 2050.085 127.120 2090.515 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 2365.085 127.120 2401.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.920 2556.325 127.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.920 -3.720 184.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 -3.720 241.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 173.405 241.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 475.765 241.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 790.765 241.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 1105.765 241.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 1420.765 241.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 1735.765 241.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 2050.765 241.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 2365.765 241.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.920 2672.605 241.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 -3.720 298.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 173.405 298.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 475.765 298.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 790.765 298.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 1105.765 298.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 1420.765 298.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 1735.765 298.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 2050.765 298.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 2365.765 298.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.920 2672.605 298.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 -3.720 355.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 173.405 355.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 475.765 355.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 790.765 355.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 1105.765 355.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 1420.765 355.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 1735.765 355.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 2050.765 355.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 2365.765 355.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.920 2672.605 355.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 -3.720 412.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 173.405 412.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 477.540 412.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 792.540 412.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 1107.540 412.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 1422.540 412.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 1737.540 412.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 2052.540 412.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 2367.540 412.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.920 2682.540 412.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 465.920 -3.720 469.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 -3.720 526.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 173.405 526.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 475.765 526.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 790.765 526.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 1105.765 526.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 1420.765 526.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 1735.765 526.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 2050.765 526.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 2365.765 526.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 522.920 2672.605 526.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 -3.720 583.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 173.405 583.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 475.765 583.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 790.765 583.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 1105.765 583.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 1420.765 583.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 1735.765 583.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 2050.765 583.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 2365.765 583.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 579.920 2672.605 583.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 -3.720 640.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 173.405 640.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 475.765 640.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 790.765 640.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 1105.765 640.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 1420.765 640.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 1735.765 640.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 2050.765 640.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 2365.765 640.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.920 2672.605 640.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 -3.720 697.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 173.405 697.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 477.540 697.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 792.540 697.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 1107.540 697.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 1422.540 697.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 1737.540 697.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 2052.540 697.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 2367.540 697.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.920 2682.540 697.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.920 -3.720 754.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 -3.720 811.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 173.405 811.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 475.765 811.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 790.765 811.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 1105.765 811.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 1420.765 811.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 1735.765 811.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 2050.765 811.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 2365.765 811.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 807.920 2672.605 811.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 -3.720 868.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 173.405 868.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 475.765 868.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 790.765 868.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 1105.765 868.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 1420.765 868.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 1735.765 868.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 2050.765 868.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 2365.765 868.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 864.920 2672.605 868.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 -3.720 925.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 173.405 925.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 475.765 925.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 790.765 925.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 1105.765 925.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 1420.765 925.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 1735.765 925.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 2050.765 925.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 2365.765 925.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.920 2672.605 925.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 -3.720 982.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 173.405 982.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 477.540 982.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 792.540 982.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 1107.540 982.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 1422.540 982.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 1737.540 982.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 2052.540 982.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 2367.540 982.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 978.920 2682.540 982.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.920 -3.720 1039.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 -3.720 1096.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 173.405 1096.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 475.765 1096.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 790.765 1096.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 1105.765 1096.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 1420.765 1096.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 1735.765 1096.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 2050.765 1096.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 2365.765 1096.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1092.920 2672.605 1096.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 -3.720 1153.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 173.405 1153.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 475.765 1153.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 790.765 1153.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 1105.765 1153.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 1420.765 1153.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 1735.765 1153.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 2050.765 1153.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 2365.765 1153.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1149.920 2672.605 1153.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 -3.720 1210.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 173.405 1210.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 475.765 1210.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 790.765 1210.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 1105.765 1210.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 1420.765 1210.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 1735.765 1210.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 2050.765 1210.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 2365.765 1210.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1206.920 2672.605 1210.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 -3.720 1267.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 173.405 1267.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 477.540 1267.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 792.540 1267.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 1107.540 1267.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 1422.540 1267.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 1737.540 1267.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 2052.540 1267.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 2367.540 1267.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.920 2682.540 1267.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1320.920 -3.720 1324.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 -3.720 1381.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 173.405 1381.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 475.765 1381.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 790.765 1381.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 1105.765 1381.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 1420.765 1381.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 1735.765 1381.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 2050.765 1381.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 2365.765 1381.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.920 2672.605 1381.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 -3.720 1438.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 173.405 1438.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 475.765 1438.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 790.765 1438.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 1105.765 1438.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 1420.765 1438.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 1735.765 1438.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 2050.765 1438.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 2365.765 1438.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1434.920 2672.605 1438.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 -3.720 1495.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 173.405 1495.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 475.765 1495.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 790.765 1495.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 1105.765 1495.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 1420.765 1495.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 1735.765 1495.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 2050.765 1495.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 2365.765 1495.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1491.920 2672.605 1495.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 -3.720 1552.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 173.405 1552.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 477.540 1552.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 792.540 1552.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 1107.540 1552.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 1422.540 1552.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 1737.540 1552.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 2052.540 1552.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 2367.540 1552.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.920 2682.540 1552.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1605.920 -3.720 1609.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 -3.720 1666.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 173.405 1666.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 475.765 1666.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 790.765 1666.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 1105.765 1666.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 1420.765 1666.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 1735.765 1666.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 2050.765 1666.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 2365.765 1666.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1662.920 2672.605 1666.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 -3.720 1723.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 173.405 1723.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 475.765 1723.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 790.765 1723.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 1105.765 1723.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 1420.765 1723.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 1735.765 1723.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 2050.765 1723.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 2365.765 1723.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.920 2672.605 1723.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 -3.720 1780.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 173.405 1780.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 475.765 1780.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 790.765 1780.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 1105.765 1780.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 1420.765 1780.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 1735.765 1780.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 2050.765 1780.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 2365.765 1780.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1776.920 2672.605 1780.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 -3.720 1837.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 173.405 1837.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 477.540 1837.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 792.540 1837.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 1107.540 1837.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 1422.540 1837.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 1737.540 1837.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 2052.540 1837.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 2367.540 1837.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1833.920 2682.540 1837.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1890.920 -3.720 1894.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 -3.720 1951.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 173.405 1951.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 475.765 1951.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 790.765 1951.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 1105.765 1951.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 1420.765 1951.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 1735.765 1951.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 2050.765 1951.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 2365.765 1951.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.920 2672.605 1951.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 -3.720 2008.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 173.405 2008.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 475.765 2008.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 790.765 2008.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 1105.765 2008.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 1420.765 2008.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 1735.765 2008.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 2050.765 2008.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 2365.765 2008.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.920 2672.605 2008.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 -3.720 2065.120 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 173.405 2065.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 475.765 2065.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 790.765 2065.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 1105.765 2065.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 1420.765 2065.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 1735.765 2065.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 2050.765 2065.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 2365.765 2065.120 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.920 2672.605 2065.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 -3.720 2122.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 173.405 2122.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 477.540 2122.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 792.540 2122.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 1107.540 2122.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 1422.540 2122.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 1737.540 2122.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 2052.540 2122.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 2367.540 2122.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2118.920 2682.540 2122.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.920 -3.720 2179.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 -3.720 2236.120 47.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 172.045 2236.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 475.765 2236.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 790.765 2236.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 1105.765 2236.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 1420.765 2236.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 1735.765 2236.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 2050.765 2236.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 2365.765 2236.120 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.920 2656.285 2236.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 -3.720 2293.120 47.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 172.045 2293.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 475.765 2293.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 790.765 2293.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 1105.765 2293.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 1420.765 2293.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 1735.765 2293.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 2050.765 2293.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 2365.765 2293.120 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.920 2656.285 2293.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 -3.720 2350.120 47.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 172.045 2350.120 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 475.765 2350.120 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 790.765 2350.120 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 1105.765 2350.120 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 1420.765 2350.120 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 1735.765 2350.120 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 2050.765 2350.120 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 2365.765 2350.120 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2346.920 2656.285 2350.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 -3.720 2407.120 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 162.940 2407.120 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 477.540 2407.120 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 792.540 2407.120 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 1107.540 2407.120 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 1422.540 2407.120 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 1737.540 2407.120 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 2052.540 2407.120 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 2367.540 2407.120 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.920 2682.540 2407.120 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2460.920 -3.720 2464.120 2718.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 25.680 2487.560 28.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 78.180 2487.560 81.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 130.680 2487.560 133.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 183.180 2487.560 186.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 235.680 2487.560 238.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 288.180 2487.560 291.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 340.680 2487.560 343.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 393.180 2487.560 396.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 445.680 2487.560 448.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 498.180 2487.560 501.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 550.680 2487.560 553.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 603.180 2487.560 606.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 655.680 2487.560 658.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 708.180 2487.560 711.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 760.680 2487.560 763.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 813.180 2487.560 816.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 865.680 2487.560 868.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 918.180 2487.560 921.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 970.680 2487.560 973.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1023.180 2487.560 1026.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1075.680 2487.560 1078.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1128.180 2487.560 1131.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1180.680 2487.560 1183.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1233.180 2487.560 1236.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1285.680 2487.560 1288.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1338.180 2487.560 1341.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1390.680 2487.560 1393.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1443.180 2487.560 1446.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1495.680 2487.560 1498.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1548.180 2487.560 1551.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1600.680 2487.560 1603.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1653.180 2487.560 1656.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1705.680 2487.560 1708.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1758.180 2487.560 1761.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1810.680 2487.560 1813.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1863.180 2487.560 1866.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1915.680 2487.560 1918.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1968.180 2487.560 1971.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2020.680 2487.560 2023.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2073.180 2487.560 2076.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2125.680 2487.560 2128.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2178.180 2487.560 2181.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2230.680 2487.560 2233.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2283.180 2487.560 2286.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2335.680 2487.560 2338.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2388.180 2487.560 2391.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2440.680 2487.560 2443.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2493.180 2487.560 2496.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2545.680 2487.560 2548.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2598.180 2487.560 2601.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2650.680 2487.560 2653.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -5.960 3.080 -1.160 2711.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.960 3.080 2480.760 7.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.960 2706.680 2480.760 2711.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.960 3.080 2480.760 2711.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.120 -3.720 8.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.120 -3.720 65.320 45.715 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.120 174.765 65.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 -3.720 122.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 174.765 122.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 477.540 122.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 792.540 122.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 1107.540 122.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 1422.540 122.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 1737.540 122.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 2052.540 122.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 2367.540 122.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.120 2682.540 122.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 176.120 -3.720 179.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 -3.720 236.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 173.405 236.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 477.540 236.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 792.540 236.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 1107.540 236.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 1422.540 236.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 1737.540 236.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 2052.540 236.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 2367.540 236.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.120 2682.540 236.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 -3.720 293.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 173.405 293.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 475.765 293.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 790.765 293.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 1105.765 293.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 1420.765 293.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 1735.765 293.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 2050.765 293.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 2365.765 293.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 290.120 2672.605 293.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 -3.720 350.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 173.405 350.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 475.765 350.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 790.765 350.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 1105.765 350.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 1420.765 350.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 1735.765 350.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 2050.765 350.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 2365.765 350.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 347.120 2672.605 350.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 -3.720 407.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 173.405 407.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 475.765 407.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 790.765 407.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 1105.765 407.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 1420.765 407.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 1735.765 407.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 2050.765 407.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 2365.765 407.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 2672.605 407.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.120 -3.720 464.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 -3.720 521.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 173.405 521.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 477.540 521.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 792.540 521.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 1107.540 521.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 1422.540 521.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 1737.540 521.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 2052.540 521.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 2367.540 521.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.120 2682.540 521.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 -3.720 578.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 173.405 578.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 475.765 578.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 790.765 578.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 1105.765 578.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 1420.765 578.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 1735.765 578.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 2050.765 578.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 2365.765 578.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.120 2672.605 578.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 -3.720 635.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 173.405 635.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 475.765 635.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 790.765 635.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 1105.765 635.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 1420.765 635.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 1735.765 635.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 2050.765 635.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 2365.765 635.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.120 2672.605 635.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 -3.720 692.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 173.405 692.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 475.765 692.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 790.765 692.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 1105.765 692.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 1420.765 692.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 1735.765 692.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 2050.765 692.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 2365.765 692.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 689.120 2672.605 692.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.120 -3.720 749.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 -3.720 806.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 173.405 806.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 477.540 806.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 792.540 806.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 1107.540 806.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 1422.540 806.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 1737.540 806.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 2052.540 806.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 2367.540 806.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.120 2682.540 806.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 -3.720 863.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 173.405 863.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 475.765 863.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 790.765 863.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 1105.765 863.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 1420.765 863.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 1735.765 863.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 2050.765 863.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 2365.765 863.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 860.120 2672.605 863.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 -3.720 920.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 173.405 920.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 475.765 920.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 790.765 920.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 1105.765 920.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 1420.765 920.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 1735.765 920.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 2050.765 920.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 2365.765 920.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.120 2672.605 920.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 -3.720 977.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 173.405 977.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 475.765 977.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 790.765 977.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 1105.765 977.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 1420.765 977.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 1735.765 977.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 2050.765 977.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 2365.765 977.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.120 2672.605 977.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1031.120 -3.720 1034.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 -3.720 1091.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 173.405 1091.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 477.540 1091.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 792.540 1091.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 1107.540 1091.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 1422.540 1091.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 1737.540 1091.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 2052.540 1091.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 2367.540 1091.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.120 2682.540 1091.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 -3.720 1148.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 173.405 1148.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 475.765 1148.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 790.765 1148.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 1105.765 1148.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 1420.765 1148.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 1735.765 1148.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 2050.765 1148.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 2365.765 1148.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1145.120 2672.605 1148.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 -3.720 1205.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 173.405 1205.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 475.765 1205.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 790.765 1205.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 1105.765 1205.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 1420.765 1205.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 1735.765 1205.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 2050.765 1205.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 2365.765 1205.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1202.120 2672.605 1205.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 -3.720 1262.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 173.405 1262.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 475.765 1262.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 790.765 1262.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 1105.765 1262.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 1420.765 1262.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 1735.765 1262.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 2050.765 1262.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 2365.765 1262.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1259.120 2672.605 1262.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1316.120 -3.720 1319.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 -3.720 1376.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 173.405 1376.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 477.540 1376.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 792.540 1376.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 1107.540 1376.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 1422.540 1376.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 1737.540 1376.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 2052.540 1376.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 2367.540 1376.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.120 2682.540 1376.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 -3.720 1433.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 173.405 1433.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 475.765 1433.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 790.765 1433.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 1105.765 1433.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 1420.765 1433.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 1735.765 1433.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 2050.765 1433.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 2365.765 1433.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1430.120 2672.605 1433.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 -3.720 1490.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 173.405 1490.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 475.765 1490.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 790.765 1490.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 1105.765 1490.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 1420.765 1490.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 1735.765 1490.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 2050.765 1490.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 2365.765 1490.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.120 2672.605 1490.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 -3.720 1547.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 173.405 1547.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 475.765 1547.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 790.765 1547.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 1105.765 1547.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 1420.765 1547.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 1735.765 1547.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 2050.765 1547.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 2365.765 1547.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.120 2672.605 1547.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1601.120 -3.720 1604.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 -3.720 1661.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 173.405 1661.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 477.540 1661.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 792.540 1661.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 1107.540 1661.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 1422.540 1661.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 1737.540 1661.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 2052.540 1661.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 2367.540 1661.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.120 2682.540 1661.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 -3.720 1718.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 173.405 1718.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 475.765 1718.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 790.765 1718.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 1105.765 1718.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 1420.765 1718.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 1735.765 1718.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 2050.765 1718.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 2365.765 1718.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1715.120 2672.605 1718.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 -3.720 1775.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 173.405 1775.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 475.765 1775.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 790.765 1775.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 1105.765 1775.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 1420.765 1775.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 1735.765 1775.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 2050.765 1775.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 2365.765 1775.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1772.120 2672.605 1775.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 -3.720 1832.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 173.405 1832.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 475.765 1832.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 790.765 1832.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 1105.765 1832.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 1420.765 1832.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 1735.765 1832.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 2050.765 1832.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 2365.765 1832.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.120 2672.605 1832.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1886.120 -3.720 1889.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 -3.720 1946.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 173.405 1946.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 477.540 1946.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 792.540 1946.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 1107.540 1946.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 1422.540 1946.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 1737.540 1946.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 2052.540 1946.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 2367.540 1946.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.120 2682.540 1946.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 -3.720 2003.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 173.405 2003.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 475.765 2003.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 790.765 2003.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 1105.765 2003.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 1420.765 2003.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 1735.765 2003.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 2050.765 2003.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 2365.765 2003.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.120 2672.605 2003.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 -3.720 2060.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 173.405 2060.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 475.765 2060.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 790.765 2060.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 1105.765 2060.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 1420.765 2060.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 1735.765 2060.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 2050.765 2060.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 2365.765 2060.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2057.120 2672.605 2060.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 -3.720 2117.320 45.035 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 173.405 2117.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 475.765 2117.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 790.765 2117.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 1105.765 2117.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 1420.765 2117.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 1735.765 2117.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 2050.765 2117.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 2365.765 2117.320 2402.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.120 2672.605 2117.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.120 -3.720 2174.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 -3.720 2231.320 30.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 172.045 2231.320 195.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 477.540 2231.320 510.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 792.540 2231.320 825.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 1107.540 2231.320 1140.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 1422.540 2231.320 1455.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 1737.540 2231.320 1770.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 2052.540 2231.320 2085.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 2367.540 2231.320 2400.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 2228.120 2682.540 2231.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 -3.720 2288.320 47.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 172.045 2288.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 475.765 2288.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 790.765 2288.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 1105.765 2288.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 1420.765 2288.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 1735.765 2288.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 2050.765 2288.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 2365.765 2288.320 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2285.120 2656.285 2288.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 -3.720 2345.320 47.755 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 172.045 2345.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 475.765 2345.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 790.765 2345.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 1105.765 2345.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 1420.765 2345.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 1735.765 2345.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 2050.765 2345.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 2365.765 2345.320 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2342.120 2656.285 2345.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 -3.720 2402.320 197.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 475.765 2402.320 512.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 790.765 2402.320 827.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 1105.765 2402.320 1142.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 1420.765 2402.320 1457.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 1735.765 2402.320 1772.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 2050.765 2402.320 2087.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 2365.765 2402.320 2402.115 ;
    END
    PORT
      LAYER met4 ;
        RECT 2399.120 2656.285 2402.320 2718.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 2456.120 -3.720 2459.320 2718.280 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 19.280 2487.560 22.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 71.780 2487.560 74.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 124.280 2487.560 127.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 176.780 2487.560 179.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 229.280 2487.560 232.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 281.780 2487.560 284.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 334.280 2487.560 337.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 386.780 2487.560 389.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 439.280 2487.560 442.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 491.780 2487.560 494.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 544.280 2487.560 547.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 596.780 2487.560 599.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 649.280 2487.560 652.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 701.780 2487.560 704.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 754.280 2487.560 757.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 806.780 2487.560 809.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 859.280 2487.560 862.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 911.780 2487.560 914.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 964.280 2487.560 967.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1016.780 2487.560 1019.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1069.280 2487.560 1072.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1121.780 2487.560 1124.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1174.280 2487.560 1177.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1226.780 2487.560 1229.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1279.280 2487.560 1282.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1331.780 2487.560 1334.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1384.280 2487.560 1387.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1436.780 2487.560 1439.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1489.280 2487.560 1492.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1541.780 2487.560 1544.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1594.280 2487.560 1597.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1646.780 2487.560 1649.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1699.280 2487.560 1702.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1751.780 2487.560 1754.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1804.280 2487.560 1807.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1856.780 2487.560 1859.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1909.280 2487.560 1912.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 1961.780 2487.560 1964.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2014.280 2487.560 2017.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2066.780 2487.560 2069.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2119.280 2487.560 2122.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2171.780 2487.560 2174.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2224.280 2487.560 2227.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2276.780 2487.560 2279.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2329.280 2487.560 2332.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2381.780 2487.560 2384.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2434.280 2487.560 2437.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2486.780 2487.560 2489.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2539.280 2487.560 2542.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2591.780 2487.560 2594.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2644.280 2487.560 2647.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.760 2696.780 2487.560 2699.980 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 2711.000 298.910 2715.000 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END clk
  PIN gfpga_pad_io_soc_dir[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 2711.000 78.110 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[0]
  PIN gfpga_pad_io_soc_dir[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END gfpga_pad_io_soc_dir[100]
  PIN gfpga_pad_io_soc_dir[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END gfpga_pad_io_soc_dir[101]
  PIN gfpga_pad_io_soc_dir[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END gfpga_pad_io_soc_dir[102]
  PIN gfpga_pad_io_soc_dir[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END gfpga_pad_io_soc_dir[103]
  PIN gfpga_pad_io_soc_dir[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END gfpga_pad_io_soc_dir[104]
  PIN gfpga_pad_io_soc_dir[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END gfpga_pad_io_soc_dir[105]
  PIN gfpga_pad_io_soc_dir[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END gfpga_pad_io_soc_dir[106]
  PIN gfpga_pad_io_soc_dir[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END gfpga_pad_io_soc_dir[107]
  PIN gfpga_pad_io_soc_dir[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END gfpga_pad_io_soc_dir[108]
  PIN gfpga_pad_io_soc_dir[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END gfpga_pad_io_soc_dir[109]
  PIN gfpga_pad_io_soc_dir[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 2711.000 784.670 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[10]
  PIN gfpga_pad_io_soc_dir[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END gfpga_pad_io_soc_dir[110]
  PIN gfpga_pad_io_soc_dir[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END gfpga_pad_io_soc_dir[111]
  PIN gfpga_pad_io_soc_dir[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END gfpga_pad_io_soc_dir[112]
  PIN gfpga_pad_io_soc_dir[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END gfpga_pad_io_soc_dir[113]
  PIN gfpga_pad_io_soc_dir[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1628.640 4.000 1629.240 ;
    END
  END gfpga_pad_io_soc_dir[114]
  PIN gfpga_pad_io_soc_dir[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END gfpga_pad_io_soc_dir[115]
  PIN gfpga_pad_io_soc_dir[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.840 4.000 1792.440 ;
    END
  END gfpga_pad_io_soc_dir[116]
  PIN gfpga_pad_io_soc_dir[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1873.440 4.000 1874.040 ;
    END
  END gfpga_pad_io_soc_dir[117]
  PIN gfpga_pad_io_soc_dir[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1955.040 4.000 1955.640 ;
    END
  END gfpga_pad_io_soc_dir[118]
  PIN gfpga_pad_io_soc_dir[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2036.640 4.000 2037.240 ;
    END
  END gfpga_pad_io_soc_dir[119]
  PIN gfpga_pad_io_soc_dir[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 2711.000 850.910 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[11]
  PIN gfpga_pad_io_soc_dir[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 4.000 2118.840 ;
    END
  END gfpga_pad_io_soc_dir[120]
  PIN gfpga_pad_io_soc_dir[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2199.840 4.000 2200.440 ;
    END
  END gfpga_pad_io_soc_dir[121]
  PIN gfpga_pad_io_soc_dir[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2281.440 4.000 2282.040 ;
    END
  END gfpga_pad_io_soc_dir[122]
  PIN gfpga_pad_io_soc_dir[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2363.040 4.000 2363.640 ;
    END
  END gfpga_pad_io_soc_dir[123]
  PIN gfpga_pad_io_soc_dir[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2444.640 4.000 2445.240 ;
    END
  END gfpga_pad_io_soc_dir[124]
  PIN gfpga_pad_io_soc_dir[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2526.240 4.000 2526.840 ;
    END
  END gfpga_pad_io_soc_dir[125]
  PIN gfpga_pad_io_soc_dir[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2607.840 4.000 2608.440 ;
    END
  END gfpga_pad_io_soc_dir[126]
  PIN gfpga_pad_io_soc_dir[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2689.440 4.000 2690.040 ;
    END
  END gfpga_pad_io_soc_dir[127]
  PIN gfpga_pad_io_soc_dir[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.870 2711.000 917.150 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[12]
  PIN gfpga_pad_io_soc_dir[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 2711.000 983.390 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[13]
  PIN gfpga_pad_io_soc_dir[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 2711.000 1049.630 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[14]
  PIN gfpga_pad_io_soc_dir[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.590 2711.000 1115.870 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[15]
  PIN gfpga_pad_io_soc_dir[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 2711.000 1182.110 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[16]
  PIN gfpga_pad_io_soc_dir[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.070 2711.000 1248.350 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[17]
  PIN gfpga_pad_io_soc_dir[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 2711.000 1314.590 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[18]
  PIN gfpga_pad_io_soc_dir[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 2711.000 1380.830 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[19]
  PIN gfpga_pad_io_soc_dir[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 2711.000 144.350 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[1]
  PIN gfpga_pad_io_soc_dir[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.790 2711.000 1447.070 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[20]
  PIN gfpga_pad_io_soc_dir[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.030 2711.000 1513.310 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[21]
  PIN gfpga_pad_io_soc_dir[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 2711.000 1579.550 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[22]
  PIN gfpga_pad_io_soc_dir[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 2711.000 1645.790 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[23]
  PIN gfpga_pad_io_soc_dir[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.750 2711.000 1712.030 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[24]
  PIN gfpga_pad_io_soc_dir[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.990 2711.000 1778.270 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[25]
  PIN gfpga_pad_io_soc_dir[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.230 2711.000 1844.510 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[26]
  PIN gfpga_pad_io_soc_dir[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.470 2711.000 1910.750 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[27]
  PIN gfpga_pad_io_soc_dir[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.710 2711.000 1976.990 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[28]
  PIN gfpga_pad_io_soc_dir[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.950 2711.000 2043.230 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[29]
  PIN gfpga_pad_io_soc_dir[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 2711.000 210.590 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[2]
  PIN gfpga_pad_io_soc_dir[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.190 2711.000 2109.470 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[30]
  PIN gfpga_pad_io_soc_dir[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.430 2711.000 2175.710 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[31]
  PIN gfpga_pad_io_soc_dir[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.670 2711.000 2241.950 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[32]
  PIN gfpga_pad_io_soc_dir[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.910 2711.000 2308.190 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[33]
  PIN gfpga_pad_io_soc_dir[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.150 2711.000 2374.430 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[34]
  PIN gfpga_pad_io_soc_dir[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.390 2711.000 2440.670 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[35]
  PIN gfpga_pad_io_soc_dir[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2590.160 2475.000 2590.760 ;
    END
  END gfpga_pad_io_soc_dir[36]
  PIN gfpga_pad_io_soc_dir[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2510.600 2475.000 2511.200 ;
    END
  END gfpga_pad_io_soc_dir[37]
  PIN gfpga_pad_io_soc_dir[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2431.040 2475.000 2431.640 ;
    END
  END gfpga_pad_io_soc_dir[38]
  PIN gfpga_pad_io_soc_dir[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2351.480 2475.000 2352.080 ;
    END
  END gfpga_pad_io_soc_dir[39]
  PIN gfpga_pad_io_soc_dir[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 2711.000 276.830 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[3]
  PIN gfpga_pad_io_soc_dir[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2271.920 2475.000 2272.520 ;
    END
  END gfpga_pad_io_soc_dir[40]
  PIN gfpga_pad_io_soc_dir[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2192.360 2475.000 2192.960 ;
    END
  END gfpga_pad_io_soc_dir[41]
  PIN gfpga_pad_io_soc_dir[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2112.800 2475.000 2113.400 ;
    END
  END gfpga_pad_io_soc_dir[42]
  PIN gfpga_pad_io_soc_dir[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2033.240 2475.000 2033.840 ;
    END
  END gfpga_pad_io_soc_dir[43]
  PIN gfpga_pad_io_soc_dir[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1953.680 2475.000 1954.280 ;
    END
  END gfpga_pad_io_soc_dir[44]
  PIN gfpga_pad_io_soc_dir[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1874.120 2475.000 1874.720 ;
    END
  END gfpga_pad_io_soc_dir[45]
  PIN gfpga_pad_io_soc_dir[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1794.560 2475.000 1795.160 ;
    END
  END gfpga_pad_io_soc_dir[46]
  PIN gfpga_pad_io_soc_dir[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1715.000 2475.000 1715.600 ;
    END
  END gfpga_pad_io_soc_dir[47]
  PIN gfpga_pad_io_soc_dir[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1635.440 2475.000 1636.040 ;
    END
  END gfpga_pad_io_soc_dir[48]
  PIN gfpga_pad_io_soc_dir[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1555.880 2475.000 1556.480 ;
    END
  END gfpga_pad_io_soc_dir[49]
  PIN gfpga_pad_io_soc_dir[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 2711.000 387.230 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[4]
  PIN gfpga_pad_io_soc_dir[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1476.320 2475.000 1476.920 ;
    END
  END gfpga_pad_io_soc_dir[50]
  PIN gfpga_pad_io_soc_dir[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1396.760 2475.000 1397.360 ;
    END
  END gfpga_pad_io_soc_dir[51]
  PIN gfpga_pad_io_soc_dir[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1317.200 2475.000 1317.800 ;
    END
  END gfpga_pad_io_soc_dir[52]
  PIN gfpga_pad_io_soc_dir[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1237.640 2475.000 1238.240 ;
    END
  END gfpga_pad_io_soc_dir[53]
  PIN gfpga_pad_io_soc_dir[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1105.040 2475.000 1105.640 ;
    END
  END gfpga_pad_io_soc_dir[54]
  PIN gfpga_pad_io_soc_dir[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1025.480 2475.000 1026.080 ;
    END
  END gfpga_pad_io_soc_dir[55]
  PIN gfpga_pad_io_soc_dir[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 945.920 2475.000 946.520 ;
    END
  END gfpga_pad_io_soc_dir[56]
  PIN gfpga_pad_io_soc_dir[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 866.360 2475.000 866.960 ;
    END
  END gfpga_pad_io_soc_dir[57]
  PIN gfpga_pad_io_soc_dir[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 786.800 2475.000 787.400 ;
    END
  END gfpga_pad_io_soc_dir[58]
  PIN gfpga_pad_io_soc_dir[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 707.240 2475.000 707.840 ;
    END
  END gfpga_pad_io_soc_dir[59]
  PIN gfpga_pad_io_soc_dir[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 2711.000 453.470 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[5]
  PIN gfpga_pad_io_soc_dir[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 627.680 2475.000 628.280 ;
    END
  END gfpga_pad_io_soc_dir[60]
  PIN gfpga_pad_io_soc_dir[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 548.120 2475.000 548.720 ;
    END
  END gfpga_pad_io_soc_dir[61]
  PIN gfpga_pad_io_soc_dir[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 468.560 2475.000 469.160 ;
    END
  END gfpga_pad_io_soc_dir[62]
  PIN gfpga_pad_io_soc_dir[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 389.000 2475.000 389.600 ;
    END
  END gfpga_pad_io_soc_dir[63]
  PIN gfpga_pad_io_soc_dir[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 309.440 2475.000 310.040 ;
    END
  END gfpga_pad_io_soc_dir[64]
  PIN gfpga_pad_io_soc_dir[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 229.880 2475.000 230.480 ;
    END
  END gfpga_pad_io_soc_dir[65]
  PIN gfpga_pad_io_soc_dir[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 150.320 2475.000 150.920 ;
    END
  END gfpga_pad_io_soc_dir[66]
  PIN gfpga_pad_io_soc_dir[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 70.760 2475.000 71.360 ;
    END
  END gfpga_pad_io_soc_dir[67]
  PIN gfpga_pad_io_soc_dir[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.230 0.000 2396.510 4.000 ;
    END
  END gfpga_pad_io_soc_dir[68]
  PIN gfpga_pad_io_soc_dir[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.290 0.000 2309.570 4.000 ;
    END
  END gfpga_pad_io_soc_dir[69]
  PIN gfpga_pad_io_soc_dir[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 2711.000 519.710 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[6]
  PIN gfpga_pad_io_soc_dir[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.350 0.000 2222.630 4.000 ;
    END
  END gfpga_pad_io_soc_dir[70]
  PIN gfpga_pad_io_soc_dir[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.410 0.000 2135.690 4.000 ;
    END
  END gfpga_pad_io_soc_dir[71]
  PIN gfpga_pad_io_soc_dir[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.470 0.000 2048.750 4.000 ;
    END
  END gfpga_pad_io_soc_dir[72]
  PIN gfpga_pad_io_soc_dir[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.530 0.000 1961.810 4.000 ;
    END
  END gfpga_pad_io_soc_dir[73]
  PIN gfpga_pad_io_soc_dir[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 0.000 1874.870 4.000 ;
    END
  END gfpga_pad_io_soc_dir[74]
  PIN gfpga_pad_io_soc_dir[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.650 0.000 1787.930 4.000 ;
    END
  END gfpga_pad_io_soc_dir[75]
  PIN gfpga_pad_io_soc_dir[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.710 0.000 1700.990 4.000 ;
    END
  END gfpga_pad_io_soc_dir[76]
  PIN gfpga_pad_io_soc_dir[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.770 0.000 1614.050 4.000 ;
    END
  END gfpga_pad_io_soc_dir[77]
  PIN gfpga_pad_io_soc_dir[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 0.000 1527.110 4.000 ;
    END
  END gfpga_pad_io_soc_dir[78]
  PIN gfpga_pad_io_soc_dir[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END gfpga_pad_io_soc_dir[79]
  PIN gfpga_pad_io_soc_dir[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 2711.000 585.950 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[7]
  PIN gfpga_pad_io_soc_dir[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END gfpga_pad_io_soc_dir[80]
  PIN gfpga_pad_io_soc_dir[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END gfpga_pad_io_soc_dir[81]
  PIN gfpga_pad_io_soc_dir[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.070 0.000 1179.350 4.000 ;
    END
  END gfpga_pad_io_soc_dir[82]
  PIN gfpga_pad_io_soc_dir[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END gfpga_pad_io_soc_dir[83]
  PIN gfpga_pad_io_soc_dir[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END gfpga_pad_io_soc_dir[84]
  PIN gfpga_pad_io_soc_dir[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 4.000 ;
    END
  END gfpga_pad_io_soc_dir[85]
  PIN gfpga_pad_io_soc_dir[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END gfpga_pad_io_soc_dir[86]
  PIN gfpga_pad_io_soc_dir[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END gfpga_pad_io_soc_dir[87]
  PIN gfpga_pad_io_soc_dir[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END gfpga_pad_io_soc_dir[88]
  PIN gfpga_pad_io_soc_dir[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END gfpga_pad_io_soc_dir[89]
  PIN gfpga_pad_io_soc_dir[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 2711.000 652.190 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[8]
  PIN gfpga_pad_io_soc_dir[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END gfpga_pad_io_soc_dir[90]
  PIN gfpga_pad_io_soc_dir[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END gfpga_pad_io_soc_dir[91]
  PIN gfpga_pad_io_soc_dir[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END gfpga_pad_io_soc_dir[92]
  PIN gfpga_pad_io_soc_dir[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END gfpga_pad_io_soc_dir[93]
  PIN gfpga_pad_io_soc_dir[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END gfpga_pad_io_soc_dir[94]
  PIN gfpga_pad_io_soc_dir[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END gfpga_pad_io_soc_dir[95]
  PIN gfpga_pad_io_soc_dir[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END gfpga_pad_io_soc_dir[96]
  PIN gfpga_pad_io_soc_dir[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END gfpga_pad_io_soc_dir[97]
  PIN gfpga_pad_io_soc_dir[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END gfpga_pad_io_soc_dir[98]
  PIN gfpga_pad_io_soc_dir[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END gfpga_pad_io_soc_dir[99]
  PIN gfpga_pad_io_soc_dir[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 2711.000 718.430 2715.000 ;
    END
  END gfpga_pad_io_soc_dir[9]
  PIN gfpga_pad_io_soc_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 2711.000 33.950 2715.000 ;
    END
  END gfpga_pad_io_soc_in[0]
  PIN gfpga_pad_io_soc_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END gfpga_pad_io_soc_in[100]
  PIN gfpga_pad_io_soc_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END gfpga_pad_io_soc_in[101]
  PIN gfpga_pad_io_soc_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END gfpga_pad_io_soc_in[102]
  PIN gfpga_pad_io_soc_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END gfpga_pad_io_soc_in[103]
  PIN gfpga_pad_io_soc_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END gfpga_pad_io_soc_in[104]
  PIN gfpga_pad_io_soc_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END gfpga_pad_io_soc_in[105]
  PIN gfpga_pad_io_soc_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END gfpga_pad_io_soc_in[106]
  PIN gfpga_pad_io_soc_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END gfpga_pad_io_soc_in[107]
  PIN gfpga_pad_io_soc_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END gfpga_pad_io_soc_in[108]
  PIN gfpga_pad_io_soc_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END gfpga_pad_io_soc_in[109]
  PIN gfpga_pad_io_soc_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 2711.000 740.510 2715.000 ;
    END
  END gfpga_pad_io_soc_in[10]
  PIN gfpga_pad_io_soc_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1220.640 4.000 1221.240 ;
    END
  END gfpga_pad_io_soc_in[110]
  PIN gfpga_pad_io_soc_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END gfpga_pad_io_soc_in[111]
  PIN gfpga_pad_io_soc_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.040 4.000 1411.640 ;
    END
  END gfpga_pad_io_soc_in[112]
  PIN gfpga_pad_io_soc_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END gfpga_pad_io_soc_in[113]
  PIN gfpga_pad_io_soc_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.240 4.000 1574.840 ;
    END
  END gfpga_pad_io_soc_in[114]
  PIN gfpga_pad_io_soc_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END gfpga_pad_io_soc_in[115]
  PIN gfpga_pad_io_soc_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1737.440 4.000 1738.040 ;
    END
  END gfpga_pad_io_soc_in[116]
  PIN gfpga_pad_io_soc_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1819.040 4.000 1819.640 ;
    END
  END gfpga_pad_io_soc_in[117]
  PIN gfpga_pad_io_soc_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1900.640 4.000 1901.240 ;
    END
  END gfpga_pad_io_soc_in[118]
  PIN gfpga_pad_io_soc_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1982.240 4.000 1982.840 ;
    END
  END gfpga_pad_io_soc_in[119]
  PIN gfpga_pad_io_soc_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 2711.000 806.750 2715.000 ;
    END
  END gfpga_pad_io_soc_in[11]
  PIN gfpga_pad_io_soc_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2063.840 4.000 2064.440 ;
    END
  END gfpga_pad_io_soc_in[120]
  PIN gfpga_pad_io_soc_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2145.440 4.000 2146.040 ;
    END
  END gfpga_pad_io_soc_in[121]
  PIN gfpga_pad_io_soc_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2227.040 4.000 2227.640 ;
    END
  END gfpga_pad_io_soc_in[122]
  PIN gfpga_pad_io_soc_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2308.640 4.000 2309.240 ;
    END
  END gfpga_pad_io_soc_in[123]
  PIN gfpga_pad_io_soc_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2390.240 4.000 2390.840 ;
    END
  END gfpga_pad_io_soc_in[124]
  PIN gfpga_pad_io_soc_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2471.840 4.000 2472.440 ;
    END
  END gfpga_pad_io_soc_in[125]
  PIN gfpga_pad_io_soc_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2553.440 4.000 2554.040 ;
    END
  END gfpga_pad_io_soc_in[126]
  PIN gfpga_pad_io_soc_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2635.040 4.000 2635.640 ;
    END
  END gfpga_pad_io_soc_in[127]
  PIN gfpga_pad_io_soc_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 2711.000 872.990 2715.000 ;
    END
  END gfpga_pad_io_soc_in[12]
  PIN gfpga_pad_io_soc_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 2711.000 939.230 2715.000 ;
    END
  END gfpga_pad_io_soc_in[13]
  PIN gfpga_pad_io_soc_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 2711.000 1005.470 2715.000 ;
    END
  END gfpga_pad_io_soc_in[14]
  PIN gfpga_pad_io_soc_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 2711.000 1071.710 2715.000 ;
    END
  END gfpga_pad_io_soc_in[15]
  PIN gfpga_pad_io_soc_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 2711.000 1137.950 2715.000 ;
    END
  END gfpga_pad_io_soc_in[16]
  PIN gfpga_pad_io_soc_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.910 2711.000 1204.190 2715.000 ;
    END
  END gfpga_pad_io_soc_in[17]
  PIN gfpga_pad_io_soc_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.150 2711.000 1270.430 2715.000 ;
    END
  END gfpga_pad_io_soc_in[18]
  PIN gfpga_pad_io_soc_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.390 2711.000 1336.670 2715.000 ;
    END
  END gfpga_pad_io_soc_in[19]
  PIN gfpga_pad_io_soc_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 2711.000 100.190 2715.000 ;
    END
  END gfpga_pad_io_soc_in[1]
  PIN gfpga_pad_io_soc_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 2711.000 1402.910 2715.000 ;
    END
  END gfpga_pad_io_soc_in[20]
  PIN gfpga_pad_io_soc_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 2711.000 1469.150 2715.000 ;
    END
  END gfpga_pad_io_soc_in[21]
  PIN gfpga_pad_io_soc_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.110 2711.000 1535.390 2715.000 ;
    END
  END gfpga_pad_io_soc_in[22]
  PIN gfpga_pad_io_soc_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.350 2711.000 1601.630 2715.000 ;
    END
  END gfpga_pad_io_soc_in[23]
  PIN gfpga_pad_io_soc_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 2711.000 1667.870 2715.000 ;
    END
  END gfpga_pad_io_soc_in[24]
  PIN gfpga_pad_io_soc_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.830 2711.000 1734.110 2715.000 ;
    END
  END gfpga_pad_io_soc_in[25]
  PIN gfpga_pad_io_soc_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 2711.000 1800.350 2715.000 ;
    END
  END gfpga_pad_io_soc_in[26]
  PIN gfpga_pad_io_soc_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.310 2711.000 1866.590 2715.000 ;
    END
  END gfpga_pad_io_soc_in[27]
  PIN gfpga_pad_io_soc_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.550 2711.000 1932.830 2715.000 ;
    END
  END gfpga_pad_io_soc_in[28]
  PIN gfpga_pad_io_soc_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.790 2711.000 1999.070 2715.000 ;
    END
  END gfpga_pad_io_soc_in[29]
  PIN gfpga_pad_io_soc_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 2711.000 166.430 2715.000 ;
    END
  END gfpga_pad_io_soc_in[2]
  PIN gfpga_pad_io_soc_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.030 2711.000 2065.310 2715.000 ;
    END
  END gfpga_pad_io_soc_in[30]
  PIN gfpga_pad_io_soc_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.270 2711.000 2131.550 2715.000 ;
    END
  END gfpga_pad_io_soc_in[31]
  PIN gfpga_pad_io_soc_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.510 2711.000 2197.790 2715.000 ;
    END
  END gfpga_pad_io_soc_in[32]
  PIN gfpga_pad_io_soc_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.750 2711.000 2264.030 2715.000 ;
    END
  END gfpga_pad_io_soc_in[33]
  PIN gfpga_pad_io_soc_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.990 2711.000 2330.270 2715.000 ;
    END
  END gfpga_pad_io_soc_in[34]
  PIN gfpga_pad_io_soc_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.230 2711.000 2396.510 2715.000 ;
    END
  END gfpga_pad_io_soc_in[35]
  PIN gfpga_pad_io_soc_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2643.200 2475.000 2643.800 ;
    END
  END gfpga_pad_io_soc_in[36]
  PIN gfpga_pad_io_soc_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2563.640 2475.000 2564.240 ;
    END
  END gfpga_pad_io_soc_in[37]
  PIN gfpga_pad_io_soc_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2484.080 2475.000 2484.680 ;
    END
  END gfpga_pad_io_soc_in[38]
  PIN gfpga_pad_io_soc_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2404.520 2475.000 2405.120 ;
    END
  END gfpga_pad_io_soc_in[39]
  PIN gfpga_pad_io_soc_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 2711.000 232.670 2715.000 ;
    END
  END gfpga_pad_io_soc_in[3]
  PIN gfpga_pad_io_soc_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2324.960 2475.000 2325.560 ;
    END
  END gfpga_pad_io_soc_in[40]
  PIN gfpga_pad_io_soc_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2245.400 2475.000 2246.000 ;
    END
  END gfpga_pad_io_soc_in[41]
  PIN gfpga_pad_io_soc_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2165.840 2475.000 2166.440 ;
    END
  END gfpga_pad_io_soc_in[42]
  PIN gfpga_pad_io_soc_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2086.280 2475.000 2086.880 ;
    END
  END gfpga_pad_io_soc_in[43]
  PIN gfpga_pad_io_soc_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2006.720 2475.000 2007.320 ;
    END
  END gfpga_pad_io_soc_in[44]
  PIN gfpga_pad_io_soc_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1927.160 2475.000 1927.760 ;
    END
  END gfpga_pad_io_soc_in[45]
  PIN gfpga_pad_io_soc_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1847.600 2475.000 1848.200 ;
    END
  END gfpga_pad_io_soc_in[46]
  PIN gfpga_pad_io_soc_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1768.040 2475.000 1768.640 ;
    END
  END gfpga_pad_io_soc_in[47]
  PIN gfpga_pad_io_soc_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1688.480 2475.000 1689.080 ;
    END
  END gfpga_pad_io_soc_in[48]
  PIN gfpga_pad_io_soc_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1608.920 2475.000 1609.520 ;
    END
  END gfpga_pad_io_soc_in[49]
  PIN gfpga_pad_io_soc_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 2711.000 343.070 2715.000 ;
    END
  END gfpga_pad_io_soc_in[4]
  PIN gfpga_pad_io_soc_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1529.360 2475.000 1529.960 ;
    END
  END gfpga_pad_io_soc_in[50]
  PIN gfpga_pad_io_soc_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1449.800 2475.000 1450.400 ;
    END
  END gfpga_pad_io_soc_in[51]
  PIN gfpga_pad_io_soc_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1370.240 2475.000 1370.840 ;
    END
  END gfpga_pad_io_soc_in[52]
  PIN gfpga_pad_io_soc_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1290.680 2475.000 1291.280 ;
    END
  END gfpga_pad_io_soc_in[53]
  PIN gfpga_pad_io_soc_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1158.080 2475.000 1158.680 ;
    END
  END gfpga_pad_io_soc_in[54]
  PIN gfpga_pad_io_soc_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1078.520 2475.000 1079.120 ;
    END
  END gfpga_pad_io_soc_in[55]
  PIN gfpga_pad_io_soc_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 998.960 2475.000 999.560 ;
    END
  END gfpga_pad_io_soc_in[56]
  PIN gfpga_pad_io_soc_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 919.400 2475.000 920.000 ;
    END
  END gfpga_pad_io_soc_in[57]
  PIN gfpga_pad_io_soc_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 839.840 2475.000 840.440 ;
    END
  END gfpga_pad_io_soc_in[58]
  PIN gfpga_pad_io_soc_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 760.280 2475.000 760.880 ;
    END
  END gfpga_pad_io_soc_in[59]
  PIN gfpga_pad_io_soc_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 2711.000 409.310 2715.000 ;
    END
  END gfpga_pad_io_soc_in[5]
  PIN gfpga_pad_io_soc_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 680.720 2475.000 681.320 ;
    END
  END gfpga_pad_io_soc_in[60]
  PIN gfpga_pad_io_soc_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 601.160 2475.000 601.760 ;
    END
  END gfpga_pad_io_soc_in[61]
  PIN gfpga_pad_io_soc_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 521.600 2475.000 522.200 ;
    END
  END gfpga_pad_io_soc_in[62]
  PIN gfpga_pad_io_soc_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 442.040 2475.000 442.640 ;
    END
  END gfpga_pad_io_soc_in[63]
  PIN gfpga_pad_io_soc_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 362.480 2475.000 363.080 ;
    END
  END gfpga_pad_io_soc_in[64]
  PIN gfpga_pad_io_soc_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 282.920 2475.000 283.520 ;
    END
  END gfpga_pad_io_soc_in[65]
  PIN gfpga_pad_io_soc_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 203.360 2475.000 203.960 ;
    END
  END gfpga_pad_io_soc_in[66]
  PIN gfpga_pad_io_soc_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 123.800 2475.000 124.400 ;
    END
  END gfpga_pad_io_soc_in[67]
  PIN gfpga_pad_io_soc_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.190 0.000 2454.470 4.000 ;
    END
  END gfpga_pad_io_soc_in[68]
  PIN gfpga_pad_io_soc_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.250 0.000 2367.530 4.000 ;
    END
  END gfpga_pad_io_soc_in[69]
  PIN gfpga_pad_io_soc_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 2711.000 475.550 2715.000 ;
    END
  END gfpga_pad_io_soc_in[6]
  PIN gfpga_pad_io_soc_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.310 0.000 2280.590 4.000 ;
    END
  END gfpga_pad_io_soc_in[70]
  PIN gfpga_pad_io_soc_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.370 0.000 2193.650 4.000 ;
    END
  END gfpga_pad_io_soc_in[71]
  PIN gfpga_pad_io_soc_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.430 0.000 2106.710 4.000 ;
    END
  END gfpga_pad_io_soc_in[72]
  PIN gfpga_pad_io_soc_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.490 0.000 2019.770 4.000 ;
    END
  END gfpga_pad_io_soc_in[73]
  PIN gfpga_pad_io_soc_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.550 0.000 1932.830 4.000 ;
    END
  END gfpga_pad_io_soc_in[74]
  PIN gfpga_pad_io_soc_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 0.000 1845.890 4.000 ;
    END
  END gfpga_pad_io_soc_in[75]
  PIN gfpga_pad_io_soc_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.670 0.000 1758.950 4.000 ;
    END
  END gfpga_pad_io_soc_in[76]
  PIN gfpga_pad_io_soc_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.730 0.000 1672.010 4.000 ;
    END
  END gfpga_pad_io_soc_in[77]
  PIN gfpga_pad_io_soc_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 0.000 1585.070 4.000 ;
    END
  END gfpga_pad_io_soc_in[78]
  PIN gfpga_pad_io_soc_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.850 0.000 1498.130 4.000 ;
    END
  END gfpga_pad_io_soc_in[79]
  PIN gfpga_pad_io_soc_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 2711.000 541.790 2715.000 ;
    END
  END gfpga_pad_io_soc_in[7]
  PIN gfpga_pad_io_soc_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 0.000 1411.190 4.000 ;
    END
  END gfpga_pad_io_soc_in[80]
  PIN gfpga_pad_io_soc_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END gfpga_pad_io_soc_in[81]
  PIN gfpga_pad_io_soc_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 0.000 1237.310 4.000 ;
    END
  END gfpga_pad_io_soc_in[82]
  PIN gfpga_pad_io_soc_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END gfpga_pad_io_soc_in[83]
  PIN gfpga_pad_io_soc_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.150 0.000 1063.430 4.000 ;
    END
  END gfpga_pad_io_soc_in[84]
  PIN gfpga_pad_io_soc_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END gfpga_pad_io_soc_in[85]
  PIN gfpga_pad_io_soc_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 0.000 889.550 4.000 ;
    END
  END gfpga_pad_io_soc_in[86]
  PIN gfpga_pad_io_soc_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END gfpga_pad_io_soc_in[87]
  PIN gfpga_pad_io_soc_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END gfpga_pad_io_soc_in[88]
  PIN gfpga_pad_io_soc_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END gfpga_pad_io_soc_in[89]
  PIN gfpga_pad_io_soc_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 2711.000 608.030 2715.000 ;
    END
  END gfpga_pad_io_soc_in[8]
  PIN gfpga_pad_io_soc_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END gfpga_pad_io_soc_in[90]
  PIN gfpga_pad_io_soc_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END gfpga_pad_io_soc_in[91]
  PIN gfpga_pad_io_soc_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END gfpga_pad_io_soc_in[92]
  PIN gfpga_pad_io_soc_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END gfpga_pad_io_soc_in[93]
  PIN gfpga_pad_io_soc_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END gfpga_pad_io_soc_in[94]
  PIN gfpga_pad_io_soc_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END gfpga_pad_io_soc_in[95]
  PIN gfpga_pad_io_soc_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END gfpga_pad_io_soc_in[96]
  PIN gfpga_pad_io_soc_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END gfpga_pad_io_soc_in[97]
  PIN gfpga_pad_io_soc_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END gfpga_pad_io_soc_in[98]
  PIN gfpga_pad_io_soc_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END gfpga_pad_io_soc_in[99]
  PIN gfpga_pad_io_soc_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 2711.000 674.270 2715.000 ;
    END
  END gfpga_pad_io_soc_in[9]
  PIN gfpga_pad_io_soc_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 2711.000 56.030 2715.000 ;
    END
  END gfpga_pad_io_soc_out[0]
  PIN gfpga_pad_io_soc_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END gfpga_pad_io_soc_out[100]
  PIN gfpga_pad_io_soc_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END gfpga_pad_io_soc_out[101]
  PIN gfpga_pad_io_soc_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END gfpga_pad_io_soc_out[102]
  PIN gfpga_pad_io_soc_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END gfpga_pad_io_soc_out[103]
  PIN gfpga_pad_io_soc_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END gfpga_pad_io_soc_out[104]
  PIN gfpga_pad_io_soc_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END gfpga_pad_io_soc_out[105]
  PIN gfpga_pad_io_soc_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END gfpga_pad_io_soc_out[106]
  PIN gfpga_pad_io_soc_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END gfpga_pad_io_soc_out[107]
  PIN gfpga_pad_io_soc_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END gfpga_pad_io_soc_out[108]
  PIN gfpga_pad_io_soc_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END gfpga_pad_io_soc_out[109]
  PIN gfpga_pad_io_soc_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 2711.000 762.590 2715.000 ;
    END
  END gfpga_pad_io_soc_out[10]
  PIN gfpga_pad_io_soc_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END gfpga_pad_io_soc_out[110]
  PIN gfpga_pad_io_soc_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1356.640 4.000 1357.240 ;
    END
  END gfpga_pad_io_soc_out[111]
  PIN gfpga_pad_io_soc_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.240 4.000 1438.840 ;
    END
  END gfpga_pad_io_soc_out[112]
  PIN gfpga_pad_io_soc_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.840 4.000 1520.440 ;
    END
  END gfpga_pad_io_soc_out[113]
  PIN gfpga_pad_io_soc_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END gfpga_pad_io_soc_out[114]
  PIN gfpga_pad_io_soc_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END gfpga_pad_io_soc_out[115]
  PIN gfpga_pad_io_soc_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1764.640 4.000 1765.240 ;
    END
  END gfpga_pad_io_soc_out[116]
  PIN gfpga_pad_io_soc_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1846.240 4.000 1846.840 ;
    END
  END gfpga_pad_io_soc_out[117]
  PIN gfpga_pad_io_soc_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END gfpga_pad_io_soc_out[118]
  PIN gfpga_pad_io_soc_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2009.440 4.000 2010.040 ;
    END
  END gfpga_pad_io_soc_out[119]
  PIN gfpga_pad_io_soc_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 2711.000 828.830 2715.000 ;
    END
  END gfpga_pad_io_soc_out[11]
  PIN gfpga_pad_io_soc_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2091.040 4.000 2091.640 ;
    END
  END gfpga_pad_io_soc_out[120]
  PIN gfpga_pad_io_soc_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2172.640 4.000 2173.240 ;
    END
  END gfpga_pad_io_soc_out[121]
  PIN gfpga_pad_io_soc_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2254.240 4.000 2254.840 ;
    END
  END gfpga_pad_io_soc_out[122]
  PIN gfpga_pad_io_soc_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2335.840 4.000 2336.440 ;
    END
  END gfpga_pad_io_soc_out[123]
  PIN gfpga_pad_io_soc_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2417.440 4.000 2418.040 ;
    END
  END gfpga_pad_io_soc_out[124]
  PIN gfpga_pad_io_soc_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2499.040 4.000 2499.640 ;
    END
  END gfpga_pad_io_soc_out[125]
  PIN gfpga_pad_io_soc_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2580.640 4.000 2581.240 ;
    END
  END gfpga_pad_io_soc_out[126]
  PIN gfpga_pad_io_soc_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2662.240 4.000 2662.840 ;
    END
  END gfpga_pad_io_soc_out[127]
  PIN gfpga_pad_io_soc_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 2711.000 895.070 2715.000 ;
    END
  END gfpga_pad_io_soc_out[12]
  PIN gfpga_pad_io_soc_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 2711.000 961.310 2715.000 ;
    END
  END gfpga_pad_io_soc_out[13]
  PIN gfpga_pad_io_soc_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.270 2711.000 1027.550 2715.000 ;
    END
  END gfpga_pad_io_soc_out[14]
  PIN gfpga_pad_io_soc_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.510 2711.000 1093.790 2715.000 ;
    END
  END gfpga_pad_io_soc_out[15]
  PIN gfpga_pad_io_soc_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.750 2711.000 1160.030 2715.000 ;
    END
  END gfpga_pad_io_soc_out[16]
  PIN gfpga_pad_io_soc_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.990 2711.000 1226.270 2715.000 ;
    END
  END gfpga_pad_io_soc_out[17]
  PIN gfpga_pad_io_soc_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.230 2711.000 1292.510 2715.000 ;
    END
  END gfpga_pad_io_soc_out[18]
  PIN gfpga_pad_io_soc_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.470 2711.000 1358.750 2715.000 ;
    END
  END gfpga_pad_io_soc_out[19]
  PIN gfpga_pad_io_soc_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 2711.000 122.270 2715.000 ;
    END
  END gfpga_pad_io_soc_out[1]
  PIN gfpga_pad_io_soc_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.710 2711.000 1424.990 2715.000 ;
    END
  END gfpga_pad_io_soc_out[20]
  PIN gfpga_pad_io_soc_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 2711.000 1491.230 2715.000 ;
    END
  END gfpga_pad_io_soc_out[21]
  PIN gfpga_pad_io_soc_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 2711.000 1557.470 2715.000 ;
    END
  END gfpga_pad_io_soc_out[22]
  PIN gfpga_pad_io_soc_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.430 2711.000 1623.710 2715.000 ;
    END
  END gfpga_pad_io_soc_out[23]
  PIN gfpga_pad_io_soc_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.670 2711.000 1689.950 2715.000 ;
    END
  END gfpga_pad_io_soc_out[24]
  PIN gfpga_pad_io_soc_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.910 2711.000 1756.190 2715.000 ;
    END
  END gfpga_pad_io_soc_out[25]
  PIN gfpga_pad_io_soc_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.150 2711.000 1822.430 2715.000 ;
    END
  END gfpga_pad_io_soc_out[26]
  PIN gfpga_pad_io_soc_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.390 2711.000 1888.670 2715.000 ;
    END
  END gfpga_pad_io_soc_out[27]
  PIN gfpga_pad_io_soc_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.630 2711.000 1954.910 2715.000 ;
    END
  END gfpga_pad_io_soc_out[28]
  PIN gfpga_pad_io_soc_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2020.870 2711.000 2021.150 2715.000 ;
    END
  END gfpga_pad_io_soc_out[29]
  PIN gfpga_pad_io_soc_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 2711.000 188.510 2715.000 ;
    END
  END gfpga_pad_io_soc_out[2]
  PIN gfpga_pad_io_soc_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2087.110 2711.000 2087.390 2715.000 ;
    END
  END gfpga_pad_io_soc_out[30]
  PIN gfpga_pad_io_soc_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.350 2711.000 2153.630 2715.000 ;
    END
  END gfpga_pad_io_soc_out[31]
  PIN gfpga_pad_io_soc_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.590 2711.000 2219.870 2715.000 ;
    END
  END gfpga_pad_io_soc_out[32]
  PIN gfpga_pad_io_soc_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2285.830 2711.000 2286.110 2715.000 ;
    END
  END gfpga_pad_io_soc_out[33]
  PIN gfpga_pad_io_soc_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.070 2711.000 2352.350 2715.000 ;
    END
  END gfpga_pad_io_soc_out[34]
  PIN gfpga_pad_io_soc_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2418.310 2711.000 2418.590 2715.000 ;
    END
  END gfpga_pad_io_soc_out[35]
  PIN gfpga_pad_io_soc_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2616.680 2475.000 2617.280 ;
    END
  END gfpga_pad_io_soc_out[36]
  PIN gfpga_pad_io_soc_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2537.120 2475.000 2537.720 ;
    END
  END gfpga_pad_io_soc_out[37]
  PIN gfpga_pad_io_soc_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2457.560 2475.000 2458.160 ;
    END
  END gfpga_pad_io_soc_out[38]
  PIN gfpga_pad_io_soc_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2378.000 2475.000 2378.600 ;
    END
  END gfpga_pad_io_soc_out[39]
  PIN gfpga_pad_io_soc_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 2711.000 254.750 2715.000 ;
    END
  END gfpga_pad_io_soc_out[3]
  PIN gfpga_pad_io_soc_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2298.440 2475.000 2299.040 ;
    END
  END gfpga_pad_io_soc_out[40]
  PIN gfpga_pad_io_soc_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2218.880 2475.000 2219.480 ;
    END
  END gfpga_pad_io_soc_out[41]
  PIN gfpga_pad_io_soc_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2139.320 2475.000 2139.920 ;
    END
  END gfpga_pad_io_soc_out[42]
  PIN gfpga_pad_io_soc_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2059.760 2475.000 2060.360 ;
    END
  END gfpga_pad_io_soc_out[43]
  PIN gfpga_pad_io_soc_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1980.200 2475.000 1980.800 ;
    END
  END gfpga_pad_io_soc_out[44]
  PIN gfpga_pad_io_soc_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1900.640 2475.000 1901.240 ;
    END
  END gfpga_pad_io_soc_out[45]
  PIN gfpga_pad_io_soc_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1821.080 2475.000 1821.680 ;
    END
  END gfpga_pad_io_soc_out[46]
  PIN gfpga_pad_io_soc_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1741.520 2475.000 1742.120 ;
    END
  END gfpga_pad_io_soc_out[47]
  PIN gfpga_pad_io_soc_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1661.960 2475.000 1662.560 ;
    END
  END gfpga_pad_io_soc_out[48]
  PIN gfpga_pad_io_soc_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1582.400 2475.000 1583.000 ;
    END
  END gfpga_pad_io_soc_out[49]
  PIN gfpga_pad_io_soc_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 2711.000 365.150 2715.000 ;
    END
  END gfpga_pad_io_soc_out[4]
  PIN gfpga_pad_io_soc_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1502.840 2475.000 1503.440 ;
    END
  END gfpga_pad_io_soc_out[50]
  PIN gfpga_pad_io_soc_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1423.280 2475.000 1423.880 ;
    END
  END gfpga_pad_io_soc_out[51]
  PIN gfpga_pad_io_soc_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1343.720 2475.000 1344.320 ;
    END
  END gfpga_pad_io_soc_out[52]
  PIN gfpga_pad_io_soc_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1264.160 2475.000 1264.760 ;
    END
  END gfpga_pad_io_soc_out[53]
  PIN gfpga_pad_io_soc_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1131.560 2475.000 1132.160 ;
    END
  END gfpga_pad_io_soc_out[54]
  PIN gfpga_pad_io_soc_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1052.000 2475.000 1052.600 ;
    END
  END gfpga_pad_io_soc_out[55]
  PIN gfpga_pad_io_soc_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 972.440 2475.000 973.040 ;
    END
  END gfpga_pad_io_soc_out[56]
  PIN gfpga_pad_io_soc_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 892.880 2475.000 893.480 ;
    END
  END gfpga_pad_io_soc_out[57]
  PIN gfpga_pad_io_soc_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 813.320 2475.000 813.920 ;
    END
  END gfpga_pad_io_soc_out[58]
  PIN gfpga_pad_io_soc_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 733.760 2475.000 734.360 ;
    END
  END gfpga_pad_io_soc_out[59]
  PIN gfpga_pad_io_soc_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 2711.000 431.390 2715.000 ;
    END
  END gfpga_pad_io_soc_out[5]
  PIN gfpga_pad_io_soc_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 654.200 2475.000 654.800 ;
    END
  END gfpga_pad_io_soc_out[60]
  PIN gfpga_pad_io_soc_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 574.640 2475.000 575.240 ;
    END
  END gfpga_pad_io_soc_out[61]
  PIN gfpga_pad_io_soc_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 495.080 2475.000 495.680 ;
    END
  END gfpga_pad_io_soc_out[62]
  PIN gfpga_pad_io_soc_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 415.520 2475.000 416.120 ;
    END
  END gfpga_pad_io_soc_out[63]
  PIN gfpga_pad_io_soc_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 335.960 2475.000 336.560 ;
    END
  END gfpga_pad_io_soc_out[64]
  PIN gfpga_pad_io_soc_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 256.400 2475.000 257.000 ;
    END
  END gfpga_pad_io_soc_out[65]
  PIN gfpga_pad_io_soc_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 176.840 2475.000 177.440 ;
    END
  END gfpga_pad_io_soc_out[66]
  PIN gfpga_pad_io_soc_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 97.280 2475.000 97.880 ;
    END
  END gfpga_pad_io_soc_out[67]
  PIN gfpga_pad_io_soc_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.210 0.000 2425.490 4.000 ;
    END
  END gfpga_pad_io_soc_out[68]
  PIN gfpga_pad_io_soc_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.270 0.000 2338.550 4.000 ;
    END
  END gfpga_pad_io_soc_out[69]
  PIN gfpga_pad_io_soc_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 2711.000 497.630 2715.000 ;
    END
  END gfpga_pad_io_soc_out[6]
  PIN gfpga_pad_io_soc_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.330 0.000 2251.610 4.000 ;
    END
  END gfpga_pad_io_soc_out[70]
  PIN gfpga_pad_io_soc_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.390 0.000 2164.670 4.000 ;
    END
  END gfpga_pad_io_soc_out[71]
  PIN gfpga_pad_io_soc_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.450 0.000 2077.730 4.000 ;
    END
  END gfpga_pad_io_soc_out[72]
  PIN gfpga_pad_io_soc_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.510 0.000 1990.790 4.000 ;
    END
  END gfpga_pad_io_soc_out[73]
  PIN gfpga_pad_io_soc_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END gfpga_pad_io_soc_out[74]
  PIN gfpga_pad_io_soc_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.630 0.000 1816.910 4.000 ;
    END
  END gfpga_pad_io_soc_out[75]
  PIN gfpga_pad_io_soc_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.690 0.000 1729.970 4.000 ;
    END
  END gfpga_pad_io_soc_out[76]
  PIN gfpga_pad_io_soc_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.750 0.000 1643.030 4.000 ;
    END
  END gfpga_pad_io_soc_out[77]
  PIN gfpga_pad_io_soc_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.810 0.000 1556.090 4.000 ;
    END
  END gfpga_pad_io_soc_out[78]
  PIN gfpga_pad_io_soc_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 0.000 1469.150 4.000 ;
    END
  END gfpga_pad_io_soc_out[79]
  PIN gfpga_pad_io_soc_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 2711.000 563.870 2715.000 ;
    END
  END gfpga_pad_io_soc_out[7]
  PIN gfpga_pad_io_soc_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 4.000 ;
    END
  END gfpga_pad_io_soc_out[80]
  PIN gfpga_pad_io_soc_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 0.000 1295.270 4.000 ;
    END
  END gfpga_pad_io_soc_out[81]
  PIN gfpga_pad_io_soc_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.050 0.000 1208.330 4.000 ;
    END
  END gfpga_pad_io_soc_out[82]
  PIN gfpga_pad_io_soc_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END gfpga_pad_io_soc_out[83]
  PIN gfpga_pad_io_soc_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END gfpga_pad_io_soc_out[84]
  PIN gfpga_pad_io_soc_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END gfpga_pad_io_soc_out[85]
  PIN gfpga_pad_io_soc_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END gfpga_pad_io_soc_out[86]
  PIN gfpga_pad_io_soc_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END gfpga_pad_io_soc_out[87]
  PIN gfpga_pad_io_soc_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END gfpga_pad_io_soc_out[88]
  PIN gfpga_pad_io_soc_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END gfpga_pad_io_soc_out[89]
  PIN gfpga_pad_io_soc_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 2711.000 630.110 2715.000 ;
    END
  END gfpga_pad_io_soc_out[8]
  PIN gfpga_pad_io_soc_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END gfpga_pad_io_soc_out[90]
  PIN gfpga_pad_io_soc_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END gfpga_pad_io_soc_out[91]
  PIN gfpga_pad_io_soc_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END gfpga_pad_io_soc_out[92]
  PIN gfpga_pad_io_soc_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END gfpga_pad_io_soc_out[93]
  PIN gfpga_pad_io_soc_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END gfpga_pad_io_soc_out[94]
  PIN gfpga_pad_io_soc_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END gfpga_pad_io_soc_out[95]
  PIN gfpga_pad_io_soc_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END gfpga_pad_io_soc_out[96]
  PIN gfpga_pad_io_soc_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END gfpga_pad_io_soc_out[97]
  PIN gfpga_pad_io_soc_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END gfpga_pad_io_soc_out[98]
  PIN gfpga_pad_io_soc_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END gfpga_pad_io_soc_out[99]
  PIN gfpga_pad_io_soc_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 2711.000 696.350 2715.000 ;
    END
  END gfpga_pad_io_soc_out[9]
  PIN isol_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 44.240 2475.000 44.840 ;
    END
  END isol_n
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END prog_clk
  PIN prog_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END prog_reset
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1184.600 2475.000 1185.200 ;
    END
  END reset
  PIN sc_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 2711.000 320.990 2715.000 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 2669.720 2475.000 2670.320 ;
    END
  END sc_tail
  PIN test_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2471.000 1211.120 2475.000 1211.720 ;
    END
  END test_enable
  OBS
      LAYER li1 ;
        RECT 1.840 10.795 2472.960 2703.765 ;
      LAYER met1 ;
        RECT 1.840 8.880 2472.960 2703.920 ;
      LAYER met2 ;
        RECT 3.310 2710.720 33.390 2711.570 ;
        RECT 34.230 2710.720 55.470 2711.570 ;
        RECT 56.310 2710.720 77.550 2711.570 ;
        RECT 78.390 2710.720 99.630 2711.570 ;
        RECT 100.470 2710.720 121.710 2711.570 ;
        RECT 122.550 2710.720 143.790 2711.570 ;
        RECT 144.630 2710.720 165.870 2711.570 ;
        RECT 166.710 2710.720 187.950 2711.570 ;
        RECT 188.790 2710.720 210.030 2711.570 ;
        RECT 210.870 2710.720 232.110 2711.570 ;
        RECT 232.950 2710.720 254.190 2711.570 ;
        RECT 255.030 2710.720 276.270 2711.570 ;
        RECT 277.110 2710.720 298.350 2711.570 ;
        RECT 299.190 2710.720 320.430 2711.570 ;
        RECT 321.270 2710.720 342.510 2711.570 ;
        RECT 343.350 2710.720 364.590 2711.570 ;
        RECT 365.430 2710.720 386.670 2711.570 ;
        RECT 387.510 2710.720 408.750 2711.570 ;
        RECT 409.590 2710.720 430.830 2711.570 ;
        RECT 431.670 2710.720 452.910 2711.570 ;
        RECT 453.750 2710.720 474.990 2711.570 ;
        RECT 475.830 2710.720 497.070 2711.570 ;
        RECT 497.910 2710.720 519.150 2711.570 ;
        RECT 519.990 2710.720 541.230 2711.570 ;
        RECT 542.070 2710.720 563.310 2711.570 ;
        RECT 564.150 2710.720 585.390 2711.570 ;
        RECT 586.230 2710.720 607.470 2711.570 ;
        RECT 608.310 2710.720 629.550 2711.570 ;
        RECT 630.390 2710.720 651.630 2711.570 ;
        RECT 652.470 2710.720 673.710 2711.570 ;
        RECT 674.550 2710.720 695.790 2711.570 ;
        RECT 696.630 2710.720 717.870 2711.570 ;
        RECT 718.710 2710.720 739.950 2711.570 ;
        RECT 740.790 2710.720 762.030 2711.570 ;
        RECT 762.870 2710.720 784.110 2711.570 ;
        RECT 784.950 2710.720 806.190 2711.570 ;
        RECT 807.030 2710.720 828.270 2711.570 ;
        RECT 829.110 2710.720 850.350 2711.570 ;
        RECT 851.190 2710.720 872.430 2711.570 ;
        RECT 873.270 2710.720 894.510 2711.570 ;
        RECT 895.350 2710.720 916.590 2711.570 ;
        RECT 917.430 2710.720 938.670 2711.570 ;
        RECT 939.510 2710.720 960.750 2711.570 ;
        RECT 961.590 2710.720 982.830 2711.570 ;
        RECT 983.670 2710.720 1004.910 2711.570 ;
        RECT 1005.750 2710.720 1026.990 2711.570 ;
        RECT 1027.830 2710.720 1049.070 2711.570 ;
        RECT 1049.910 2710.720 1071.150 2711.570 ;
        RECT 1071.990 2710.720 1093.230 2711.570 ;
        RECT 1094.070 2710.720 1115.310 2711.570 ;
        RECT 1116.150 2710.720 1137.390 2711.570 ;
        RECT 1138.230 2710.720 1159.470 2711.570 ;
        RECT 1160.310 2710.720 1181.550 2711.570 ;
        RECT 1182.390 2710.720 1203.630 2711.570 ;
        RECT 1204.470 2710.720 1225.710 2711.570 ;
        RECT 1226.550 2710.720 1247.790 2711.570 ;
        RECT 1248.630 2710.720 1269.870 2711.570 ;
        RECT 1270.710 2710.720 1291.950 2711.570 ;
        RECT 1292.790 2710.720 1314.030 2711.570 ;
        RECT 1314.870 2710.720 1336.110 2711.570 ;
        RECT 1336.950 2710.720 1358.190 2711.570 ;
        RECT 1359.030 2710.720 1380.270 2711.570 ;
        RECT 1381.110 2710.720 1402.350 2711.570 ;
        RECT 1403.190 2710.720 1424.430 2711.570 ;
        RECT 1425.270 2710.720 1446.510 2711.570 ;
        RECT 1447.350 2710.720 1468.590 2711.570 ;
        RECT 1469.430 2710.720 1490.670 2711.570 ;
        RECT 1491.510 2710.720 1512.750 2711.570 ;
        RECT 1513.590 2710.720 1534.830 2711.570 ;
        RECT 1535.670 2710.720 1556.910 2711.570 ;
        RECT 1557.750 2710.720 1578.990 2711.570 ;
        RECT 1579.830 2710.720 1601.070 2711.570 ;
        RECT 1601.910 2710.720 1623.150 2711.570 ;
        RECT 1623.990 2710.720 1645.230 2711.570 ;
        RECT 1646.070 2710.720 1667.310 2711.570 ;
        RECT 1668.150 2710.720 1689.390 2711.570 ;
        RECT 1690.230 2710.720 1711.470 2711.570 ;
        RECT 1712.310 2710.720 1733.550 2711.570 ;
        RECT 1734.390 2710.720 1755.630 2711.570 ;
        RECT 1756.470 2710.720 1777.710 2711.570 ;
        RECT 1778.550 2710.720 1799.790 2711.570 ;
        RECT 1800.630 2710.720 1821.870 2711.570 ;
        RECT 1822.710 2710.720 1843.950 2711.570 ;
        RECT 1844.790 2710.720 1866.030 2711.570 ;
        RECT 1866.870 2710.720 1888.110 2711.570 ;
        RECT 1888.950 2710.720 1910.190 2711.570 ;
        RECT 1911.030 2710.720 1932.270 2711.570 ;
        RECT 1933.110 2710.720 1954.350 2711.570 ;
        RECT 1955.190 2710.720 1976.430 2711.570 ;
        RECT 1977.270 2710.720 1998.510 2711.570 ;
        RECT 1999.350 2710.720 2020.590 2711.570 ;
        RECT 2021.430 2710.720 2042.670 2711.570 ;
        RECT 2043.510 2710.720 2064.750 2711.570 ;
        RECT 2065.590 2710.720 2086.830 2711.570 ;
        RECT 2087.670 2710.720 2108.910 2711.570 ;
        RECT 2109.750 2710.720 2130.990 2711.570 ;
        RECT 2131.830 2710.720 2153.070 2711.570 ;
        RECT 2153.910 2710.720 2175.150 2711.570 ;
        RECT 2175.990 2710.720 2197.230 2711.570 ;
        RECT 2198.070 2710.720 2219.310 2711.570 ;
        RECT 2220.150 2710.720 2241.390 2711.570 ;
        RECT 2242.230 2710.720 2263.470 2711.570 ;
        RECT 2264.310 2710.720 2285.550 2711.570 ;
        RECT 2286.390 2710.720 2307.630 2711.570 ;
        RECT 2308.470 2710.720 2329.710 2711.570 ;
        RECT 2330.550 2710.720 2351.790 2711.570 ;
        RECT 2352.630 2710.720 2373.870 2711.570 ;
        RECT 2374.710 2710.720 2395.950 2711.570 ;
        RECT 2396.790 2710.720 2418.030 2711.570 ;
        RECT 2418.870 2710.720 2440.110 2711.570 ;
        RECT 2440.950 2710.720 2471.020 2711.570 ;
        RECT 3.310 4.280 2471.020 2710.720 ;
        RECT 3.310 3.670 19.590 4.280 ;
        RECT 20.430 3.670 48.570 4.280 ;
        RECT 49.410 3.670 77.550 4.280 ;
        RECT 78.390 3.670 106.530 4.280 ;
        RECT 107.370 3.670 135.510 4.280 ;
        RECT 136.350 3.670 164.490 4.280 ;
        RECT 165.330 3.670 193.470 4.280 ;
        RECT 194.310 3.670 222.450 4.280 ;
        RECT 223.290 3.670 251.430 4.280 ;
        RECT 252.270 3.670 280.410 4.280 ;
        RECT 281.250 3.670 309.390 4.280 ;
        RECT 310.230 3.670 338.370 4.280 ;
        RECT 339.210 3.670 367.350 4.280 ;
        RECT 368.190 3.670 396.330 4.280 ;
        RECT 397.170 3.670 425.310 4.280 ;
        RECT 426.150 3.670 454.290 4.280 ;
        RECT 455.130 3.670 483.270 4.280 ;
        RECT 484.110 3.670 512.250 4.280 ;
        RECT 513.090 3.670 541.230 4.280 ;
        RECT 542.070 3.670 570.210 4.280 ;
        RECT 571.050 3.670 599.190 4.280 ;
        RECT 600.030 3.670 628.170 4.280 ;
        RECT 629.010 3.670 657.150 4.280 ;
        RECT 657.990 3.670 686.130 4.280 ;
        RECT 686.970 3.670 715.110 4.280 ;
        RECT 715.950 3.670 744.090 4.280 ;
        RECT 744.930 3.670 773.070 4.280 ;
        RECT 773.910 3.670 802.050 4.280 ;
        RECT 802.890 3.670 831.030 4.280 ;
        RECT 831.870 3.670 860.010 4.280 ;
        RECT 860.850 3.670 888.990 4.280 ;
        RECT 889.830 3.670 917.970 4.280 ;
        RECT 918.810 3.670 946.950 4.280 ;
        RECT 947.790 3.670 975.930 4.280 ;
        RECT 976.770 3.670 1004.910 4.280 ;
        RECT 1005.750 3.670 1033.890 4.280 ;
        RECT 1034.730 3.670 1062.870 4.280 ;
        RECT 1063.710 3.670 1091.850 4.280 ;
        RECT 1092.690 3.670 1120.830 4.280 ;
        RECT 1121.670 3.670 1149.810 4.280 ;
        RECT 1150.650 3.670 1178.790 4.280 ;
        RECT 1179.630 3.670 1207.770 4.280 ;
        RECT 1208.610 3.670 1236.750 4.280 ;
        RECT 1237.590 3.670 1265.730 4.280 ;
        RECT 1266.570 3.670 1294.710 4.280 ;
        RECT 1295.550 3.670 1323.690 4.280 ;
        RECT 1324.530 3.670 1352.670 4.280 ;
        RECT 1353.510 3.670 1381.650 4.280 ;
        RECT 1382.490 3.670 1410.630 4.280 ;
        RECT 1411.470 3.670 1439.610 4.280 ;
        RECT 1440.450 3.670 1468.590 4.280 ;
        RECT 1469.430 3.670 1497.570 4.280 ;
        RECT 1498.410 3.670 1526.550 4.280 ;
        RECT 1527.390 3.670 1555.530 4.280 ;
        RECT 1556.370 3.670 1584.510 4.280 ;
        RECT 1585.350 3.670 1613.490 4.280 ;
        RECT 1614.330 3.670 1642.470 4.280 ;
        RECT 1643.310 3.670 1671.450 4.280 ;
        RECT 1672.290 3.670 1700.430 4.280 ;
        RECT 1701.270 3.670 1729.410 4.280 ;
        RECT 1730.250 3.670 1758.390 4.280 ;
        RECT 1759.230 3.670 1787.370 4.280 ;
        RECT 1788.210 3.670 1816.350 4.280 ;
        RECT 1817.190 3.670 1845.330 4.280 ;
        RECT 1846.170 3.670 1874.310 4.280 ;
        RECT 1875.150 3.670 1903.290 4.280 ;
        RECT 1904.130 3.670 1932.270 4.280 ;
        RECT 1933.110 3.670 1961.250 4.280 ;
        RECT 1962.090 3.670 1990.230 4.280 ;
        RECT 1991.070 3.670 2019.210 4.280 ;
        RECT 2020.050 3.670 2048.190 4.280 ;
        RECT 2049.030 3.670 2077.170 4.280 ;
        RECT 2078.010 3.670 2106.150 4.280 ;
        RECT 2106.990 3.670 2135.130 4.280 ;
        RECT 2135.970 3.670 2164.110 4.280 ;
        RECT 2164.950 3.670 2193.090 4.280 ;
        RECT 2193.930 3.670 2222.070 4.280 ;
        RECT 2222.910 3.670 2251.050 4.280 ;
        RECT 2251.890 3.670 2280.030 4.280 ;
        RECT 2280.870 3.670 2309.010 4.280 ;
        RECT 2309.850 3.670 2337.990 4.280 ;
        RECT 2338.830 3.670 2366.970 4.280 ;
        RECT 2367.810 3.670 2395.950 4.280 ;
        RECT 2396.790 3.670 2424.930 4.280 ;
        RECT 2425.770 3.670 2453.910 4.280 ;
        RECT 2454.750 3.670 2471.020 4.280 ;
      LAYER met3 ;
        RECT 3.285 2690.440 2471.000 2703.845 ;
        RECT 4.400 2689.040 2471.000 2690.440 ;
        RECT 3.285 2670.720 2471.000 2689.040 ;
        RECT 3.285 2669.320 2470.600 2670.720 ;
        RECT 3.285 2663.240 2471.000 2669.320 ;
        RECT 4.400 2661.840 2471.000 2663.240 ;
        RECT 3.285 2644.200 2471.000 2661.840 ;
        RECT 3.285 2642.800 2470.600 2644.200 ;
        RECT 3.285 2636.040 2471.000 2642.800 ;
        RECT 4.400 2634.640 2471.000 2636.040 ;
        RECT 3.285 2617.680 2471.000 2634.640 ;
        RECT 3.285 2616.280 2470.600 2617.680 ;
        RECT 3.285 2608.840 2471.000 2616.280 ;
        RECT 4.400 2607.440 2471.000 2608.840 ;
        RECT 3.285 2591.160 2471.000 2607.440 ;
        RECT 3.285 2589.760 2470.600 2591.160 ;
        RECT 3.285 2581.640 2471.000 2589.760 ;
        RECT 4.400 2580.240 2471.000 2581.640 ;
        RECT 3.285 2564.640 2471.000 2580.240 ;
        RECT 3.285 2563.240 2470.600 2564.640 ;
        RECT 3.285 2554.440 2471.000 2563.240 ;
        RECT 4.400 2553.040 2471.000 2554.440 ;
        RECT 3.285 2538.120 2471.000 2553.040 ;
        RECT 3.285 2536.720 2470.600 2538.120 ;
        RECT 3.285 2527.240 2471.000 2536.720 ;
        RECT 4.400 2525.840 2471.000 2527.240 ;
        RECT 3.285 2511.600 2471.000 2525.840 ;
        RECT 3.285 2510.200 2470.600 2511.600 ;
        RECT 3.285 2500.040 2471.000 2510.200 ;
        RECT 4.400 2498.640 2471.000 2500.040 ;
        RECT 3.285 2485.080 2471.000 2498.640 ;
        RECT 3.285 2483.680 2470.600 2485.080 ;
        RECT 3.285 2472.840 2471.000 2483.680 ;
        RECT 4.400 2471.440 2471.000 2472.840 ;
        RECT 3.285 2458.560 2471.000 2471.440 ;
        RECT 3.285 2457.160 2470.600 2458.560 ;
        RECT 3.285 2445.640 2471.000 2457.160 ;
        RECT 4.400 2444.240 2471.000 2445.640 ;
        RECT 3.285 2432.040 2471.000 2444.240 ;
        RECT 3.285 2430.640 2470.600 2432.040 ;
        RECT 3.285 2418.440 2471.000 2430.640 ;
        RECT 4.400 2417.040 2471.000 2418.440 ;
        RECT 3.285 2405.520 2471.000 2417.040 ;
        RECT 3.285 2404.120 2470.600 2405.520 ;
        RECT 3.285 2391.240 2471.000 2404.120 ;
        RECT 4.400 2389.840 2471.000 2391.240 ;
        RECT 3.285 2379.000 2471.000 2389.840 ;
        RECT 3.285 2377.600 2470.600 2379.000 ;
        RECT 3.285 2364.040 2471.000 2377.600 ;
        RECT 4.400 2362.640 2471.000 2364.040 ;
        RECT 3.285 2352.480 2471.000 2362.640 ;
        RECT 3.285 2351.080 2470.600 2352.480 ;
        RECT 3.285 2336.840 2471.000 2351.080 ;
        RECT 4.400 2335.440 2471.000 2336.840 ;
        RECT 3.285 2325.960 2471.000 2335.440 ;
        RECT 3.285 2324.560 2470.600 2325.960 ;
        RECT 3.285 2309.640 2471.000 2324.560 ;
        RECT 4.400 2308.240 2471.000 2309.640 ;
        RECT 3.285 2299.440 2471.000 2308.240 ;
        RECT 3.285 2298.040 2470.600 2299.440 ;
        RECT 3.285 2282.440 2471.000 2298.040 ;
        RECT 4.400 2281.040 2471.000 2282.440 ;
        RECT 3.285 2272.920 2471.000 2281.040 ;
        RECT 3.285 2271.520 2470.600 2272.920 ;
        RECT 3.285 2255.240 2471.000 2271.520 ;
        RECT 4.400 2253.840 2471.000 2255.240 ;
        RECT 3.285 2246.400 2471.000 2253.840 ;
        RECT 3.285 2245.000 2470.600 2246.400 ;
        RECT 3.285 2228.040 2471.000 2245.000 ;
        RECT 4.400 2226.640 2471.000 2228.040 ;
        RECT 3.285 2219.880 2471.000 2226.640 ;
        RECT 3.285 2218.480 2470.600 2219.880 ;
        RECT 3.285 2200.840 2471.000 2218.480 ;
        RECT 4.400 2199.440 2471.000 2200.840 ;
        RECT 3.285 2193.360 2471.000 2199.440 ;
        RECT 3.285 2191.960 2470.600 2193.360 ;
        RECT 3.285 2173.640 2471.000 2191.960 ;
        RECT 4.400 2172.240 2471.000 2173.640 ;
        RECT 3.285 2166.840 2471.000 2172.240 ;
        RECT 3.285 2165.440 2470.600 2166.840 ;
        RECT 3.285 2146.440 2471.000 2165.440 ;
        RECT 4.400 2145.040 2471.000 2146.440 ;
        RECT 3.285 2140.320 2471.000 2145.040 ;
        RECT 3.285 2138.920 2470.600 2140.320 ;
        RECT 3.285 2119.240 2471.000 2138.920 ;
        RECT 4.400 2117.840 2471.000 2119.240 ;
        RECT 3.285 2113.800 2471.000 2117.840 ;
        RECT 3.285 2112.400 2470.600 2113.800 ;
        RECT 3.285 2092.040 2471.000 2112.400 ;
        RECT 4.400 2090.640 2471.000 2092.040 ;
        RECT 3.285 2087.280 2471.000 2090.640 ;
        RECT 3.285 2085.880 2470.600 2087.280 ;
        RECT 3.285 2064.840 2471.000 2085.880 ;
        RECT 4.400 2063.440 2471.000 2064.840 ;
        RECT 3.285 2060.760 2471.000 2063.440 ;
        RECT 3.285 2059.360 2470.600 2060.760 ;
        RECT 3.285 2037.640 2471.000 2059.360 ;
        RECT 4.400 2036.240 2471.000 2037.640 ;
        RECT 3.285 2034.240 2471.000 2036.240 ;
        RECT 3.285 2032.840 2470.600 2034.240 ;
        RECT 3.285 2010.440 2471.000 2032.840 ;
        RECT 4.400 2009.040 2471.000 2010.440 ;
        RECT 3.285 2007.720 2471.000 2009.040 ;
        RECT 3.285 2006.320 2470.600 2007.720 ;
        RECT 3.285 1983.240 2471.000 2006.320 ;
        RECT 4.400 1981.840 2471.000 1983.240 ;
        RECT 3.285 1981.200 2471.000 1981.840 ;
        RECT 3.285 1979.800 2470.600 1981.200 ;
        RECT 3.285 1956.040 2471.000 1979.800 ;
        RECT 4.400 1954.680 2471.000 1956.040 ;
        RECT 4.400 1954.640 2470.600 1954.680 ;
        RECT 3.285 1953.280 2470.600 1954.640 ;
        RECT 3.285 1928.840 2471.000 1953.280 ;
        RECT 4.400 1928.160 2471.000 1928.840 ;
        RECT 4.400 1927.440 2470.600 1928.160 ;
        RECT 3.285 1926.760 2470.600 1927.440 ;
        RECT 3.285 1901.640 2471.000 1926.760 ;
        RECT 4.400 1900.240 2470.600 1901.640 ;
        RECT 3.285 1875.120 2471.000 1900.240 ;
        RECT 3.285 1874.440 2470.600 1875.120 ;
        RECT 4.400 1873.720 2470.600 1874.440 ;
        RECT 4.400 1873.040 2471.000 1873.720 ;
        RECT 3.285 1848.600 2471.000 1873.040 ;
        RECT 3.285 1847.240 2470.600 1848.600 ;
        RECT 4.400 1847.200 2470.600 1847.240 ;
        RECT 4.400 1845.840 2471.000 1847.200 ;
        RECT 3.285 1822.080 2471.000 1845.840 ;
        RECT 3.285 1820.680 2470.600 1822.080 ;
        RECT 3.285 1820.040 2471.000 1820.680 ;
        RECT 4.400 1818.640 2471.000 1820.040 ;
        RECT 3.285 1795.560 2471.000 1818.640 ;
        RECT 3.285 1794.160 2470.600 1795.560 ;
        RECT 3.285 1792.840 2471.000 1794.160 ;
        RECT 4.400 1791.440 2471.000 1792.840 ;
        RECT 3.285 1769.040 2471.000 1791.440 ;
        RECT 3.285 1767.640 2470.600 1769.040 ;
        RECT 3.285 1765.640 2471.000 1767.640 ;
        RECT 4.400 1764.240 2471.000 1765.640 ;
        RECT 3.285 1742.520 2471.000 1764.240 ;
        RECT 3.285 1741.120 2470.600 1742.520 ;
        RECT 3.285 1738.440 2471.000 1741.120 ;
        RECT 4.400 1737.040 2471.000 1738.440 ;
        RECT 3.285 1716.000 2471.000 1737.040 ;
        RECT 3.285 1714.600 2470.600 1716.000 ;
        RECT 3.285 1711.240 2471.000 1714.600 ;
        RECT 4.400 1709.840 2471.000 1711.240 ;
        RECT 3.285 1689.480 2471.000 1709.840 ;
        RECT 3.285 1688.080 2470.600 1689.480 ;
        RECT 3.285 1684.040 2471.000 1688.080 ;
        RECT 4.400 1682.640 2471.000 1684.040 ;
        RECT 3.285 1662.960 2471.000 1682.640 ;
        RECT 3.285 1661.560 2470.600 1662.960 ;
        RECT 3.285 1656.840 2471.000 1661.560 ;
        RECT 4.400 1655.440 2471.000 1656.840 ;
        RECT 3.285 1636.440 2471.000 1655.440 ;
        RECT 3.285 1635.040 2470.600 1636.440 ;
        RECT 3.285 1629.640 2471.000 1635.040 ;
        RECT 4.400 1628.240 2471.000 1629.640 ;
        RECT 3.285 1609.920 2471.000 1628.240 ;
        RECT 3.285 1608.520 2470.600 1609.920 ;
        RECT 3.285 1602.440 2471.000 1608.520 ;
        RECT 4.400 1601.040 2471.000 1602.440 ;
        RECT 3.285 1583.400 2471.000 1601.040 ;
        RECT 3.285 1582.000 2470.600 1583.400 ;
        RECT 3.285 1575.240 2471.000 1582.000 ;
        RECT 4.400 1573.840 2471.000 1575.240 ;
        RECT 3.285 1556.880 2471.000 1573.840 ;
        RECT 3.285 1555.480 2470.600 1556.880 ;
        RECT 3.285 1548.040 2471.000 1555.480 ;
        RECT 4.400 1546.640 2471.000 1548.040 ;
        RECT 3.285 1530.360 2471.000 1546.640 ;
        RECT 3.285 1528.960 2470.600 1530.360 ;
        RECT 3.285 1520.840 2471.000 1528.960 ;
        RECT 4.400 1519.440 2471.000 1520.840 ;
        RECT 3.285 1503.840 2471.000 1519.440 ;
        RECT 3.285 1502.440 2470.600 1503.840 ;
        RECT 3.285 1493.640 2471.000 1502.440 ;
        RECT 4.400 1492.240 2471.000 1493.640 ;
        RECT 3.285 1477.320 2471.000 1492.240 ;
        RECT 3.285 1475.920 2470.600 1477.320 ;
        RECT 3.285 1466.440 2471.000 1475.920 ;
        RECT 4.400 1465.040 2471.000 1466.440 ;
        RECT 3.285 1450.800 2471.000 1465.040 ;
        RECT 3.285 1449.400 2470.600 1450.800 ;
        RECT 3.285 1439.240 2471.000 1449.400 ;
        RECT 4.400 1437.840 2471.000 1439.240 ;
        RECT 3.285 1424.280 2471.000 1437.840 ;
        RECT 3.285 1422.880 2470.600 1424.280 ;
        RECT 3.285 1412.040 2471.000 1422.880 ;
        RECT 4.400 1410.640 2471.000 1412.040 ;
        RECT 3.285 1397.760 2471.000 1410.640 ;
        RECT 3.285 1396.360 2470.600 1397.760 ;
        RECT 3.285 1384.840 2471.000 1396.360 ;
        RECT 4.400 1383.440 2471.000 1384.840 ;
        RECT 3.285 1371.240 2471.000 1383.440 ;
        RECT 3.285 1369.840 2470.600 1371.240 ;
        RECT 3.285 1357.640 2471.000 1369.840 ;
        RECT 4.400 1356.240 2471.000 1357.640 ;
        RECT 3.285 1344.720 2471.000 1356.240 ;
        RECT 3.285 1343.320 2470.600 1344.720 ;
        RECT 3.285 1330.440 2471.000 1343.320 ;
        RECT 4.400 1329.040 2471.000 1330.440 ;
        RECT 3.285 1318.200 2471.000 1329.040 ;
        RECT 3.285 1316.800 2470.600 1318.200 ;
        RECT 3.285 1303.240 2471.000 1316.800 ;
        RECT 4.400 1301.840 2471.000 1303.240 ;
        RECT 3.285 1291.680 2471.000 1301.840 ;
        RECT 3.285 1290.280 2470.600 1291.680 ;
        RECT 3.285 1276.040 2471.000 1290.280 ;
        RECT 4.400 1274.640 2471.000 1276.040 ;
        RECT 3.285 1265.160 2471.000 1274.640 ;
        RECT 3.285 1263.760 2470.600 1265.160 ;
        RECT 3.285 1248.840 2471.000 1263.760 ;
        RECT 4.400 1247.440 2471.000 1248.840 ;
        RECT 3.285 1238.640 2471.000 1247.440 ;
        RECT 3.285 1237.240 2470.600 1238.640 ;
        RECT 3.285 1221.640 2471.000 1237.240 ;
        RECT 4.400 1220.240 2471.000 1221.640 ;
        RECT 3.285 1212.120 2471.000 1220.240 ;
        RECT 3.285 1210.720 2470.600 1212.120 ;
        RECT 3.285 1194.440 2471.000 1210.720 ;
        RECT 4.400 1193.040 2471.000 1194.440 ;
        RECT 3.285 1185.600 2471.000 1193.040 ;
        RECT 3.285 1184.200 2470.600 1185.600 ;
        RECT 3.285 1167.240 2471.000 1184.200 ;
        RECT 4.400 1165.840 2471.000 1167.240 ;
        RECT 3.285 1159.080 2471.000 1165.840 ;
        RECT 3.285 1157.680 2470.600 1159.080 ;
        RECT 3.285 1140.040 2471.000 1157.680 ;
        RECT 4.400 1138.640 2471.000 1140.040 ;
        RECT 3.285 1132.560 2471.000 1138.640 ;
        RECT 3.285 1131.160 2470.600 1132.560 ;
        RECT 3.285 1112.840 2471.000 1131.160 ;
        RECT 4.400 1111.440 2471.000 1112.840 ;
        RECT 3.285 1106.040 2471.000 1111.440 ;
        RECT 3.285 1104.640 2470.600 1106.040 ;
        RECT 3.285 1085.640 2471.000 1104.640 ;
        RECT 4.400 1084.240 2471.000 1085.640 ;
        RECT 3.285 1079.520 2471.000 1084.240 ;
        RECT 3.285 1078.120 2470.600 1079.520 ;
        RECT 3.285 1058.440 2471.000 1078.120 ;
        RECT 4.400 1057.040 2471.000 1058.440 ;
        RECT 3.285 1053.000 2471.000 1057.040 ;
        RECT 3.285 1051.600 2470.600 1053.000 ;
        RECT 3.285 1031.240 2471.000 1051.600 ;
        RECT 4.400 1029.840 2471.000 1031.240 ;
        RECT 3.285 1026.480 2471.000 1029.840 ;
        RECT 3.285 1025.080 2470.600 1026.480 ;
        RECT 3.285 1004.040 2471.000 1025.080 ;
        RECT 4.400 1002.640 2471.000 1004.040 ;
        RECT 3.285 999.960 2471.000 1002.640 ;
        RECT 3.285 998.560 2470.600 999.960 ;
        RECT 3.285 976.840 2471.000 998.560 ;
        RECT 4.400 975.440 2471.000 976.840 ;
        RECT 3.285 973.440 2471.000 975.440 ;
        RECT 3.285 972.040 2470.600 973.440 ;
        RECT 3.285 949.640 2471.000 972.040 ;
        RECT 4.400 948.240 2471.000 949.640 ;
        RECT 3.285 946.920 2471.000 948.240 ;
        RECT 3.285 945.520 2470.600 946.920 ;
        RECT 3.285 922.440 2471.000 945.520 ;
        RECT 4.400 921.040 2471.000 922.440 ;
        RECT 3.285 920.400 2471.000 921.040 ;
        RECT 3.285 919.000 2470.600 920.400 ;
        RECT 3.285 895.240 2471.000 919.000 ;
        RECT 4.400 893.880 2471.000 895.240 ;
        RECT 4.400 893.840 2470.600 893.880 ;
        RECT 3.285 892.480 2470.600 893.840 ;
        RECT 3.285 868.040 2471.000 892.480 ;
        RECT 4.400 867.360 2471.000 868.040 ;
        RECT 4.400 866.640 2470.600 867.360 ;
        RECT 3.285 865.960 2470.600 866.640 ;
        RECT 3.285 840.840 2471.000 865.960 ;
        RECT 4.400 839.440 2470.600 840.840 ;
        RECT 3.285 814.320 2471.000 839.440 ;
        RECT 3.285 813.640 2470.600 814.320 ;
        RECT 4.400 812.920 2470.600 813.640 ;
        RECT 4.400 812.240 2471.000 812.920 ;
        RECT 3.285 787.800 2471.000 812.240 ;
        RECT 3.285 786.440 2470.600 787.800 ;
        RECT 4.400 786.400 2470.600 786.440 ;
        RECT 4.400 785.040 2471.000 786.400 ;
        RECT 3.285 761.280 2471.000 785.040 ;
        RECT 3.285 759.880 2470.600 761.280 ;
        RECT 3.285 759.240 2471.000 759.880 ;
        RECT 4.400 757.840 2471.000 759.240 ;
        RECT 3.285 734.760 2471.000 757.840 ;
        RECT 3.285 733.360 2470.600 734.760 ;
        RECT 3.285 732.040 2471.000 733.360 ;
        RECT 4.400 730.640 2471.000 732.040 ;
        RECT 3.285 708.240 2471.000 730.640 ;
        RECT 3.285 706.840 2470.600 708.240 ;
        RECT 3.285 704.840 2471.000 706.840 ;
        RECT 4.400 703.440 2471.000 704.840 ;
        RECT 3.285 681.720 2471.000 703.440 ;
        RECT 3.285 680.320 2470.600 681.720 ;
        RECT 3.285 677.640 2471.000 680.320 ;
        RECT 4.400 676.240 2471.000 677.640 ;
        RECT 3.285 655.200 2471.000 676.240 ;
        RECT 3.285 653.800 2470.600 655.200 ;
        RECT 3.285 650.440 2471.000 653.800 ;
        RECT 4.400 649.040 2471.000 650.440 ;
        RECT 3.285 628.680 2471.000 649.040 ;
        RECT 3.285 627.280 2470.600 628.680 ;
        RECT 3.285 623.240 2471.000 627.280 ;
        RECT 4.400 621.840 2471.000 623.240 ;
        RECT 3.285 602.160 2471.000 621.840 ;
        RECT 3.285 600.760 2470.600 602.160 ;
        RECT 3.285 596.040 2471.000 600.760 ;
        RECT 4.400 594.640 2471.000 596.040 ;
        RECT 3.285 575.640 2471.000 594.640 ;
        RECT 3.285 574.240 2470.600 575.640 ;
        RECT 3.285 568.840 2471.000 574.240 ;
        RECT 4.400 567.440 2471.000 568.840 ;
        RECT 3.285 549.120 2471.000 567.440 ;
        RECT 3.285 547.720 2470.600 549.120 ;
        RECT 3.285 541.640 2471.000 547.720 ;
        RECT 4.400 540.240 2471.000 541.640 ;
        RECT 3.285 522.600 2471.000 540.240 ;
        RECT 3.285 521.200 2470.600 522.600 ;
        RECT 3.285 514.440 2471.000 521.200 ;
        RECT 4.400 513.040 2471.000 514.440 ;
        RECT 3.285 496.080 2471.000 513.040 ;
        RECT 3.285 494.680 2470.600 496.080 ;
        RECT 3.285 487.240 2471.000 494.680 ;
        RECT 4.400 485.840 2471.000 487.240 ;
        RECT 3.285 469.560 2471.000 485.840 ;
        RECT 3.285 468.160 2470.600 469.560 ;
        RECT 3.285 460.040 2471.000 468.160 ;
        RECT 4.400 458.640 2471.000 460.040 ;
        RECT 3.285 443.040 2471.000 458.640 ;
        RECT 3.285 441.640 2470.600 443.040 ;
        RECT 3.285 432.840 2471.000 441.640 ;
        RECT 4.400 431.440 2471.000 432.840 ;
        RECT 3.285 416.520 2471.000 431.440 ;
        RECT 3.285 415.120 2470.600 416.520 ;
        RECT 3.285 405.640 2471.000 415.120 ;
        RECT 4.400 404.240 2471.000 405.640 ;
        RECT 3.285 390.000 2471.000 404.240 ;
        RECT 3.285 388.600 2470.600 390.000 ;
        RECT 3.285 378.440 2471.000 388.600 ;
        RECT 4.400 377.040 2471.000 378.440 ;
        RECT 3.285 363.480 2471.000 377.040 ;
        RECT 3.285 362.080 2470.600 363.480 ;
        RECT 3.285 351.240 2471.000 362.080 ;
        RECT 4.400 349.840 2471.000 351.240 ;
        RECT 3.285 336.960 2471.000 349.840 ;
        RECT 3.285 335.560 2470.600 336.960 ;
        RECT 3.285 324.040 2471.000 335.560 ;
        RECT 4.400 322.640 2471.000 324.040 ;
        RECT 3.285 310.440 2471.000 322.640 ;
        RECT 3.285 309.040 2470.600 310.440 ;
        RECT 3.285 296.840 2471.000 309.040 ;
        RECT 4.400 295.440 2471.000 296.840 ;
        RECT 3.285 283.920 2471.000 295.440 ;
        RECT 3.285 282.520 2470.600 283.920 ;
        RECT 3.285 269.640 2471.000 282.520 ;
        RECT 4.400 268.240 2471.000 269.640 ;
        RECT 3.285 257.400 2471.000 268.240 ;
        RECT 3.285 256.000 2470.600 257.400 ;
        RECT 3.285 242.440 2471.000 256.000 ;
        RECT 4.400 241.040 2471.000 242.440 ;
        RECT 3.285 230.880 2471.000 241.040 ;
        RECT 3.285 229.480 2470.600 230.880 ;
        RECT 3.285 215.240 2471.000 229.480 ;
        RECT 4.400 213.840 2471.000 215.240 ;
        RECT 3.285 204.360 2471.000 213.840 ;
        RECT 3.285 202.960 2470.600 204.360 ;
        RECT 3.285 188.040 2471.000 202.960 ;
        RECT 4.400 186.640 2471.000 188.040 ;
        RECT 3.285 177.840 2471.000 186.640 ;
        RECT 3.285 176.440 2470.600 177.840 ;
        RECT 3.285 160.840 2471.000 176.440 ;
        RECT 4.400 159.440 2471.000 160.840 ;
        RECT 3.285 151.320 2471.000 159.440 ;
        RECT 3.285 149.920 2470.600 151.320 ;
        RECT 3.285 133.640 2471.000 149.920 ;
        RECT 4.400 132.240 2471.000 133.640 ;
        RECT 3.285 124.800 2471.000 132.240 ;
        RECT 3.285 123.400 2470.600 124.800 ;
        RECT 3.285 106.440 2471.000 123.400 ;
        RECT 4.400 105.040 2471.000 106.440 ;
        RECT 3.285 98.280 2471.000 105.040 ;
        RECT 3.285 96.880 2470.600 98.280 ;
        RECT 3.285 79.240 2471.000 96.880 ;
        RECT 4.400 77.840 2471.000 79.240 ;
        RECT 3.285 71.760 2471.000 77.840 ;
        RECT 3.285 70.360 2470.600 71.760 ;
        RECT 3.285 52.040 2471.000 70.360 ;
        RECT 4.400 50.640 2471.000 52.040 ;
        RECT 3.285 45.240 2471.000 50.640 ;
        RECT 3.285 43.840 2470.600 45.240 ;
        RECT 3.285 24.840 2471.000 43.840 ;
        RECT 4.400 23.440 2471.000 24.840 ;
        RECT 3.285 10.715 2471.000 23.440 ;
      LAYER met4 ;
        RECT 41.335 174.365 61.720 2672.240 ;
        RECT 65.720 2555.925 123.520 2672.240 ;
        RECT 127.520 2555.925 175.720 2672.240 ;
        RECT 65.720 2401.835 175.720 2555.925 ;
        RECT 65.720 2400.740 123.520 2401.835 ;
        RECT 65.720 2367.140 66.520 2400.740 ;
        RECT 70.520 2367.140 118.720 2400.740 ;
        RECT 122.720 2367.140 123.520 2400.740 ;
        RECT 65.720 2364.685 123.520 2367.140 ;
        RECT 127.520 2364.685 175.720 2401.835 ;
        RECT 65.720 2090.915 175.720 2364.685 ;
        RECT 65.720 2085.740 123.520 2090.915 ;
        RECT 65.720 2052.140 66.520 2085.740 ;
        RECT 70.520 2052.140 118.720 2085.740 ;
        RECT 122.720 2052.140 123.520 2085.740 ;
        RECT 65.720 2049.685 123.520 2052.140 ;
        RECT 127.520 2049.685 175.720 2090.915 ;
        RECT 65.720 1775.915 175.720 2049.685 ;
        RECT 65.720 1770.740 123.520 1775.915 ;
        RECT 65.720 1737.140 66.520 1770.740 ;
        RECT 70.520 1737.140 118.720 1770.740 ;
        RECT 122.720 1737.140 123.520 1770.740 ;
        RECT 65.720 1734.685 123.520 1737.140 ;
        RECT 127.520 1734.685 175.720 1775.915 ;
        RECT 65.720 1460.915 175.720 1734.685 ;
        RECT 65.720 1455.740 123.520 1460.915 ;
        RECT 65.720 1422.140 66.520 1455.740 ;
        RECT 70.520 1422.140 118.720 1455.740 ;
        RECT 122.720 1422.140 123.520 1455.740 ;
        RECT 65.720 1419.685 123.520 1422.140 ;
        RECT 127.520 1419.685 175.720 1460.915 ;
        RECT 65.720 1145.915 175.720 1419.685 ;
        RECT 65.720 1140.740 123.520 1145.915 ;
        RECT 65.720 1107.140 66.520 1140.740 ;
        RECT 70.520 1107.140 118.720 1140.740 ;
        RECT 122.720 1107.140 123.520 1140.740 ;
        RECT 65.720 1104.685 123.520 1107.140 ;
        RECT 127.520 1104.685 175.720 1145.915 ;
        RECT 65.720 830.915 175.720 1104.685 ;
        RECT 65.720 825.740 123.520 830.915 ;
        RECT 65.720 792.140 66.520 825.740 ;
        RECT 70.520 792.140 118.720 825.740 ;
        RECT 122.720 792.140 123.520 825.740 ;
        RECT 65.720 789.685 123.520 792.140 ;
        RECT 127.520 789.685 175.720 830.915 ;
        RECT 65.720 515.915 175.720 789.685 ;
        RECT 65.720 510.740 123.520 515.915 ;
        RECT 65.720 477.140 66.520 510.740 ;
        RECT 70.520 477.140 118.720 510.740 ;
        RECT 122.720 477.140 123.520 510.740 ;
        RECT 65.720 474.685 123.520 477.140 ;
        RECT 127.520 474.685 175.720 515.915 ;
        RECT 65.720 200.915 175.720 474.685 ;
        RECT 65.720 195.740 123.520 200.915 ;
        RECT 65.720 174.365 66.520 195.740 ;
        RECT 70.520 174.365 118.720 195.740 ;
        RECT 122.720 174.365 123.520 195.740 ;
        RECT 127.520 174.365 175.720 200.915 ;
        RECT 41.335 46.115 175.720 174.365 ;
        RECT 41.335 40.640 61.720 46.115 ;
        RECT 65.720 40.640 123.520 46.115 ;
        RECT 127.520 40.640 175.720 46.115 ;
        RECT 179.720 40.640 180.520 2672.240 ;
        RECT 184.520 2672.205 237.520 2672.240 ;
        RECT 241.520 2672.205 289.720 2672.240 ;
        RECT 293.720 2672.205 294.520 2672.240 ;
        RECT 298.520 2672.205 346.720 2672.240 ;
        RECT 350.720 2672.205 351.520 2672.240 ;
        RECT 355.520 2672.205 403.720 2672.240 ;
        RECT 407.720 2672.205 460.720 2672.240 ;
        RECT 184.520 2403.195 460.720 2672.205 ;
        RECT 184.520 2400.740 237.520 2403.195 ;
        RECT 184.520 2367.140 232.720 2400.740 ;
        RECT 236.720 2367.140 237.520 2400.740 ;
        RECT 184.520 2365.365 237.520 2367.140 ;
        RECT 241.520 2365.365 289.720 2403.195 ;
        RECT 293.720 2365.365 294.520 2403.195 ;
        RECT 298.520 2365.365 346.720 2403.195 ;
        RECT 350.720 2365.365 351.520 2403.195 ;
        RECT 355.520 2365.365 403.720 2403.195 ;
        RECT 407.720 2400.740 460.720 2403.195 ;
        RECT 407.720 2367.140 408.520 2400.740 ;
        RECT 412.520 2367.140 460.720 2400.740 ;
        RECT 407.720 2365.365 460.720 2367.140 ;
        RECT 184.520 2087.515 460.720 2365.365 ;
        RECT 184.520 2085.740 237.520 2087.515 ;
        RECT 184.520 2052.140 232.720 2085.740 ;
        RECT 236.720 2052.140 237.520 2085.740 ;
        RECT 184.520 2050.365 237.520 2052.140 ;
        RECT 241.520 2050.365 289.720 2087.515 ;
        RECT 293.720 2050.365 294.520 2087.515 ;
        RECT 298.520 2050.365 346.720 2087.515 ;
        RECT 350.720 2050.365 351.520 2087.515 ;
        RECT 355.520 2050.365 403.720 2087.515 ;
        RECT 407.720 2085.740 460.720 2087.515 ;
        RECT 407.720 2052.140 408.520 2085.740 ;
        RECT 412.520 2052.140 460.720 2085.740 ;
        RECT 407.720 2050.365 460.720 2052.140 ;
        RECT 184.520 1772.515 460.720 2050.365 ;
        RECT 184.520 1770.740 237.520 1772.515 ;
        RECT 184.520 1737.140 232.720 1770.740 ;
        RECT 236.720 1737.140 237.520 1770.740 ;
        RECT 184.520 1735.365 237.520 1737.140 ;
        RECT 241.520 1735.365 289.720 1772.515 ;
        RECT 293.720 1735.365 294.520 1772.515 ;
        RECT 298.520 1735.365 346.720 1772.515 ;
        RECT 350.720 1735.365 351.520 1772.515 ;
        RECT 355.520 1735.365 403.720 1772.515 ;
        RECT 407.720 1770.740 460.720 1772.515 ;
        RECT 407.720 1737.140 408.520 1770.740 ;
        RECT 412.520 1737.140 460.720 1770.740 ;
        RECT 407.720 1735.365 460.720 1737.140 ;
        RECT 184.520 1457.515 460.720 1735.365 ;
        RECT 184.520 1455.740 237.520 1457.515 ;
        RECT 184.520 1422.140 232.720 1455.740 ;
        RECT 236.720 1422.140 237.520 1455.740 ;
        RECT 184.520 1420.365 237.520 1422.140 ;
        RECT 241.520 1420.365 289.720 1457.515 ;
        RECT 293.720 1420.365 294.520 1457.515 ;
        RECT 298.520 1420.365 346.720 1457.515 ;
        RECT 350.720 1420.365 351.520 1457.515 ;
        RECT 355.520 1420.365 403.720 1457.515 ;
        RECT 407.720 1455.740 460.720 1457.515 ;
        RECT 407.720 1422.140 408.520 1455.740 ;
        RECT 412.520 1422.140 460.720 1455.740 ;
        RECT 407.720 1420.365 460.720 1422.140 ;
        RECT 184.520 1142.515 460.720 1420.365 ;
        RECT 184.520 1140.740 237.520 1142.515 ;
        RECT 184.520 1107.140 232.720 1140.740 ;
        RECT 236.720 1107.140 237.520 1140.740 ;
        RECT 184.520 1105.365 237.520 1107.140 ;
        RECT 241.520 1105.365 289.720 1142.515 ;
        RECT 293.720 1105.365 294.520 1142.515 ;
        RECT 298.520 1105.365 346.720 1142.515 ;
        RECT 350.720 1105.365 351.520 1142.515 ;
        RECT 355.520 1105.365 403.720 1142.515 ;
        RECT 407.720 1140.740 460.720 1142.515 ;
        RECT 407.720 1107.140 408.520 1140.740 ;
        RECT 412.520 1107.140 460.720 1140.740 ;
        RECT 407.720 1105.365 460.720 1107.140 ;
        RECT 184.520 827.515 460.720 1105.365 ;
        RECT 184.520 825.740 237.520 827.515 ;
        RECT 184.520 792.140 232.720 825.740 ;
        RECT 236.720 792.140 237.520 825.740 ;
        RECT 184.520 790.365 237.520 792.140 ;
        RECT 241.520 790.365 289.720 827.515 ;
        RECT 293.720 790.365 294.520 827.515 ;
        RECT 298.520 790.365 346.720 827.515 ;
        RECT 350.720 790.365 351.520 827.515 ;
        RECT 355.520 790.365 403.720 827.515 ;
        RECT 407.720 825.740 460.720 827.515 ;
        RECT 407.720 792.140 408.520 825.740 ;
        RECT 412.520 792.140 460.720 825.740 ;
        RECT 407.720 790.365 460.720 792.140 ;
        RECT 184.520 512.515 460.720 790.365 ;
        RECT 184.520 510.740 237.520 512.515 ;
        RECT 184.520 477.140 232.720 510.740 ;
        RECT 236.720 477.140 237.520 510.740 ;
        RECT 184.520 475.365 237.520 477.140 ;
        RECT 241.520 475.365 289.720 512.515 ;
        RECT 293.720 475.365 294.520 512.515 ;
        RECT 298.520 475.365 346.720 512.515 ;
        RECT 350.720 475.365 351.520 512.515 ;
        RECT 355.520 475.365 403.720 512.515 ;
        RECT 407.720 510.740 460.720 512.515 ;
        RECT 407.720 477.140 408.520 510.740 ;
        RECT 412.520 477.140 460.720 510.740 ;
        RECT 407.720 475.365 460.720 477.140 ;
        RECT 184.520 197.515 460.720 475.365 ;
        RECT 184.520 195.740 237.520 197.515 ;
        RECT 184.520 173.005 232.720 195.740 ;
        RECT 236.720 173.005 237.520 195.740 ;
        RECT 241.520 173.005 289.720 197.515 ;
        RECT 293.720 173.005 294.520 197.515 ;
        RECT 298.520 173.005 346.720 197.515 ;
        RECT 350.720 173.005 351.520 197.515 ;
        RECT 355.520 173.005 403.720 197.515 ;
        RECT 407.720 195.740 460.720 197.515 ;
        RECT 407.720 173.005 408.520 195.740 ;
        RECT 412.520 173.005 460.720 195.740 ;
        RECT 184.520 45.435 460.720 173.005 ;
        RECT 184.520 40.640 237.520 45.435 ;
        RECT 241.520 40.640 289.720 45.435 ;
        RECT 293.720 40.640 294.520 45.435 ;
        RECT 298.520 40.640 346.720 45.435 ;
        RECT 350.720 40.640 351.520 45.435 ;
        RECT 355.520 40.640 403.720 45.435 ;
        RECT 407.720 40.640 460.720 45.435 ;
        RECT 464.720 40.640 465.520 2672.240 ;
        RECT 469.520 2672.205 522.520 2672.240 ;
        RECT 526.520 2672.205 574.720 2672.240 ;
        RECT 578.720 2672.205 579.520 2672.240 ;
        RECT 583.520 2672.205 631.720 2672.240 ;
        RECT 635.720 2672.205 636.520 2672.240 ;
        RECT 640.520 2672.205 688.720 2672.240 ;
        RECT 692.720 2672.205 745.720 2672.240 ;
        RECT 469.520 2403.195 745.720 2672.205 ;
        RECT 469.520 2400.740 522.520 2403.195 ;
        RECT 469.520 2367.140 517.720 2400.740 ;
        RECT 521.720 2367.140 522.520 2400.740 ;
        RECT 469.520 2365.365 522.520 2367.140 ;
        RECT 526.520 2365.365 574.720 2403.195 ;
        RECT 578.720 2365.365 579.520 2403.195 ;
        RECT 583.520 2365.365 631.720 2403.195 ;
        RECT 635.720 2365.365 636.520 2403.195 ;
        RECT 640.520 2365.365 688.720 2403.195 ;
        RECT 692.720 2400.740 745.720 2403.195 ;
        RECT 692.720 2367.140 693.520 2400.740 ;
        RECT 697.520 2367.140 745.720 2400.740 ;
        RECT 692.720 2365.365 745.720 2367.140 ;
        RECT 469.520 2087.515 745.720 2365.365 ;
        RECT 469.520 2085.740 522.520 2087.515 ;
        RECT 469.520 2052.140 517.720 2085.740 ;
        RECT 521.720 2052.140 522.520 2085.740 ;
        RECT 469.520 2050.365 522.520 2052.140 ;
        RECT 526.520 2050.365 574.720 2087.515 ;
        RECT 578.720 2050.365 579.520 2087.515 ;
        RECT 583.520 2050.365 631.720 2087.515 ;
        RECT 635.720 2050.365 636.520 2087.515 ;
        RECT 640.520 2050.365 688.720 2087.515 ;
        RECT 692.720 2085.740 745.720 2087.515 ;
        RECT 692.720 2052.140 693.520 2085.740 ;
        RECT 697.520 2052.140 745.720 2085.740 ;
        RECT 692.720 2050.365 745.720 2052.140 ;
        RECT 469.520 1772.515 745.720 2050.365 ;
        RECT 469.520 1770.740 522.520 1772.515 ;
        RECT 469.520 1737.140 517.720 1770.740 ;
        RECT 521.720 1737.140 522.520 1770.740 ;
        RECT 469.520 1735.365 522.520 1737.140 ;
        RECT 526.520 1735.365 574.720 1772.515 ;
        RECT 578.720 1735.365 579.520 1772.515 ;
        RECT 583.520 1735.365 631.720 1772.515 ;
        RECT 635.720 1735.365 636.520 1772.515 ;
        RECT 640.520 1735.365 688.720 1772.515 ;
        RECT 692.720 1770.740 745.720 1772.515 ;
        RECT 692.720 1737.140 693.520 1770.740 ;
        RECT 697.520 1737.140 745.720 1770.740 ;
        RECT 692.720 1735.365 745.720 1737.140 ;
        RECT 469.520 1457.515 745.720 1735.365 ;
        RECT 469.520 1455.740 522.520 1457.515 ;
        RECT 469.520 1422.140 517.720 1455.740 ;
        RECT 521.720 1422.140 522.520 1455.740 ;
        RECT 469.520 1420.365 522.520 1422.140 ;
        RECT 526.520 1420.365 574.720 1457.515 ;
        RECT 578.720 1420.365 579.520 1457.515 ;
        RECT 583.520 1420.365 631.720 1457.515 ;
        RECT 635.720 1420.365 636.520 1457.515 ;
        RECT 640.520 1420.365 688.720 1457.515 ;
        RECT 692.720 1455.740 745.720 1457.515 ;
        RECT 692.720 1422.140 693.520 1455.740 ;
        RECT 697.520 1422.140 745.720 1455.740 ;
        RECT 692.720 1420.365 745.720 1422.140 ;
        RECT 469.520 1142.515 745.720 1420.365 ;
        RECT 469.520 1140.740 522.520 1142.515 ;
        RECT 469.520 1107.140 517.720 1140.740 ;
        RECT 521.720 1107.140 522.520 1140.740 ;
        RECT 469.520 1105.365 522.520 1107.140 ;
        RECT 526.520 1105.365 574.720 1142.515 ;
        RECT 578.720 1105.365 579.520 1142.515 ;
        RECT 583.520 1105.365 631.720 1142.515 ;
        RECT 635.720 1105.365 636.520 1142.515 ;
        RECT 640.520 1105.365 688.720 1142.515 ;
        RECT 692.720 1140.740 745.720 1142.515 ;
        RECT 692.720 1107.140 693.520 1140.740 ;
        RECT 697.520 1107.140 745.720 1140.740 ;
        RECT 692.720 1105.365 745.720 1107.140 ;
        RECT 469.520 827.515 745.720 1105.365 ;
        RECT 469.520 825.740 522.520 827.515 ;
        RECT 469.520 792.140 517.720 825.740 ;
        RECT 521.720 792.140 522.520 825.740 ;
        RECT 469.520 790.365 522.520 792.140 ;
        RECT 526.520 790.365 574.720 827.515 ;
        RECT 578.720 790.365 579.520 827.515 ;
        RECT 583.520 790.365 631.720 827.515 ;
        RECT 635.720 790.365 636.520 827.515 ;
        RECT 640.520 790.365 688.720 827.515 ;
        RECT 692.720 825.740 745.720 827.515 ;
        RECT 692.720 792.140 693.520 825.740 ;
        RECT 697.520 792.140 745.720 825.740 ;
        RECT 692.720 790.365 745.720 792.140 ;
        RECT 469.520 512.515 745.720 790.365 ;
        RECT 469.520 510.740 522.520 512.515 ;
        RECT 469.520 477.140 517.720 510.740 ;
        RECT 521.720 477.140 522.520 510.740 ;
        RECT 469.520 475.365 522.520 477.140 ;
        RECT 526.520 475.365 574.720 512.515 ;
        RECT 578.720 475.365 579.520 512.515 ;
        RECT 583.520 475.365 631.720 512.515 ;
        RECT 635.720 475.365 636.520 512.515 ;
        RECT 640.520 475.365 688.720 512.515 ;
        RECT 692.720 510.740 745.720 512.515 ;
        RECT 692.720 477.140 693.520 510.740 ;
        RECT 697.520 477.140 745.720 510.740 ;
        RECT 692.720 475.365 745.720 477.140 ;
        RECT 469.520 197.515 745.720 475.365 ;
        RECT 469.520 195.740 522.520 197.515 ;
        RECT 469.520 173.005 517.720 195.740 ;
        RECT 521.720 173.005 522.520 195.740 ;
        RECT 526.520 173.005 574.720 197.515 ;
        RECT 578.720 173.005 579.520 197.515 ;
        RECT 583.520 173.005 631.720 197.515 ;
        RECT 635.720 173.005 636.520 197.515 ;
        RECT 640.520 173.005 688.720 197.515 ;
        RECT 692.720 195.740 745.720 197.515 ;
        RECT 692.720 173.005 693.520 195.740 ;
        RECT 697.520 173.005 745.720 195.740 ;
        RECT 469.520 45.435 745.720 173.005 ;
        RECT 469.520 40.640 522.520 45.435 ;
        RECT 526.520 40.640 574.720 45.435 ;
        RECT 578.720 40.640 579.520 45.435 ;
        RECT 583.520 40.640 631.720 45.435 ;
        RECT 635.720 40.640 636.520 45.435 ;
        RECT 640.520 40.640 688.720 45.435 ;
        RECT 692.720 40.640 745.720 45.435 ;
        RECT 749.720 40.640 750.520 2672.240 ;
        RECT 754.520 2672.205 807.520 2672.240 ;
        RECT 811.520 2672.205 859.720 2672.240 ;
        RECT 863.720 2672.205 864.520 2672.240 ;
        RECT 868.520 2672.205 916.720 2672.240 ;
        RECT 920.720 2672.205 921.520 2672.240 ;
        RECT 925.520 2672.205 973.720 2672.240 ;
        RECT 977.720 2672.205 1030.720 2672.240 ;
        RECT 754.520 2403.195 1030.720 2672.205 ;
        RECT 754.520 2400.740 807.520 2403.195 ;
        RECT 754.520 2367.140 802.720 2400.740 ;
        RECT 806.720 2367.140 807.520 2400.740 ;
        RECT 754.520 2365.365 807.520 2367.140 ;
        RECT 811.520 2365.365 859.720 2403.195 ;
        RECT 863.720 2365.365 864.520 2403.195 ;
        RECT 868.520 2365.365 916.720 2403.195 ;
        RECT 920.720 2365.365 921.520 2403.195 ;
        RECT 925.520 2365.365 973.720 2403.195 ;
        RECT 977.720 2400.740 1030.720 2403.195 ;
        RECT 977.720 2367.140 978.520 2400.740 ;
        RECT 982.520 2367.140 1030.720 2400.740 ;
        RECT 977.720 2365.365 1030.720 2367.140 ;
        RECT 754.520 2087.515 1030.720 2365.365 ;
        RECT 754.520 2085.740 807.520 2087.515 ;
        RECT 754.520 2052.140 802.720 2085.740 ;
        RECT 806.720 2052.140 807.520 2085.740 ;
        RECT 754.520 2050.365 807.520 2052.140 ;
        RECT 811.520 2050.365 859.720 2087.515 ;
        RECT 863.720 2050.365 864.520 2087.515 ;
        RECT 868.520 2050.365 916.720 2087.515 ;
        RECT 920.720 2050.365 921.520 2087.515 ;
        RECT 925.520 2050.365 973.720 2087.515 ;
        RECT 977.720 2085.740 1030.720 2087.515 ;
        RECT 977.720 2052.140 978.520 2085.740 ;
        RECT 982.520 2052.140 1030.720 2085.740 ;
        RECT 977.720 2050.365 1030.720 2052.140 ;
        RECT 754.520 1772.515 1030.720 2050.365 ;
        RECT 754.520 1770.740 807.520 1772.515 ;
        RECT 754.520 1737.140 802.720 1770.740 ;
        RECT 806.720 1737.140 807.520 1770.740 ;
        RECT 754.520 1735.365 807.520 1737.140 ;
        RECT 811.520 1735.365 859.720 1772.515 ;
        RECT 863.720 1735.365 864.520 1772.515 ;
        RECT 868.520 1735.365 916.720 1772.515 ;
        RECT 920.720 1735.365 921.520 1772.515 ;
        RECT 925.520 1735.365 973.720 1772.515 ;
        RECT 977.720 1770.740 1030.720 1772.515 ;
        RECT 977.720 1737.140 978.520 1770.740 ;
        RECT 982.520 1737.140 1030.720 1770.740 ;
        RECT 977.720 1735.365 1030.720 1737.140 ;
        RECT 754.520 1457.515 1030.720 1735.365 ;
        RECT 754.520 1455.740 807.520 1457.515 ;
        RECT 754.520 1422.140 802.720 1455.740 ;
        RECT 806.720 1422.140 807.520 1455.740 ;
        RECT 754.520 1420.365 807.520 1422.140 ;
        RECT 811.520 1420.365 859.720 1457.515 ;
        RECT 863.720 1420.365 864.520 1457.515 ;
        RECT 868.520 1420.365 916.720 1457.515 ;
        RECT 920.720 1420.365 921.520 1457.515 ;
        RECT 925.520 1420.365 973.720 1457.515 ;
        RECT 977.720 1455.740 1030.720 1457.515 ;
        RECT 977.720 1422.140 978.520 1455.740 ;
        RECT 982.520 1422.140 1030.720 1455.740 ;
        RECT 977.720 1420.365 1030.720 1422.140 ;
        RECT 754.520 1142.515 1030.720 1420.365 ;
        RECT 754.520 1140.740 807.520 1142.515 ;
        RECT 754.520 1107.140 802.720 1140.740 ;
        RECT 806.720 1107.140 807.520 1140.740 ;
        RECT 754.520 1105.365 807.520 1107.140 ;
        RECT 811.520 1105.365 859.720 1142.515 ;
        RECT 863.720 1105.365 864.520 1142.515 ;
        RECT 868.520 1105.365 916.720 1142.515 ;
        RECT 920.720 1105.365 921.520 1142.515 ;
        RECT 925.520 1105.365 973.720 1142.515 ;
        RECT 977.720 1140.740 1030.720 1142.515 ;
        RECT 977.720 1107.140 978.520 1140.740 ;
        RECT 982.520 1107.140 1030.720 1140.740 ;
        RECT 977.720 1105.365 1030.720 1107.140 ;
        RECT 754.520 827.515 1030.720 1105.365 ;
        RECT 754.520 825.740 807.520 827.515 ;
        RECT 754.520 792.140 802.720 825.740 ;
        RECT 806.720 792.140 807.520 825.740 ;
        RECT 754.520 790.365 807.520 792.140 ;
        RECT 811.520 790.365 859.720 827.515 ;
        RECT 863.720 790.365 864.520 827.515 ;
        RECT 868.520 790.365 916.720 827.515 ;
        RECT 920.720 790.365 921.520 827.515 ;
        RECT 925.520 790.365 973.720 827.515 ;
        RECT 977.720 825.740 1030.720 827.515 ;
        RECT 977.720 792.140 978.520 825.740 ;
        RECT 982.520 792.140 1030.720 825.740 ;
        RECT 977.720 790.365 1030.720 792.140 ;
        RECT 754.520 512.515 1030.720 790.365 ;
        RECT 754.520 510.740 807.520 512.515 ;
        RECT 754.520 477.140 802.720 510.740 ;
        RECT 806.720 477.140 807.520 510.740 ;
        RECT 754.520 475.365 807.520 477.140 ;
        RECT 811.520 475.365 859.720 512.515 ;
        RECT 863.720 475.365 864.520 512.515 ;
        RECT 868.520 475.365 916.720 512.515 ;
        RECT 920.720 475.365 921.520 512.515 ;
        RECT 925.520 475.365 973.720 512.515 ;
        RECT 977.720 510.740 1030.720 512.515 ;
        RECT 977.720 477.140 978.520 510.740 ;
        RECT 982.520 477.140 1030.720 510.740 ;
        RECT 977.720 475.365 1030.720 477.140 ;
        RECT 754.520 197.515 1030.720 475.365 ;
        RECT 754.520 195.740 807.520 197.515 ;
        RECT 754.520 173.005 802.720 195.740 ;
        RECT 806.720 173.005 807.520 195.740 ;
        RECT 811.520 173.005 859.720 197.515 ;
        RECT 863.720 173.005 864.520 197.515 ;
        RECT 868.520 173.005 916.720 197.515 ;
        RECT 920.720 173.005 921.520 197.515 ;
        RECT 925.520 173.005 973.720 197.515 ;
        RECT 977.720 195.740 1030.720 197.515 ;
        RECT 977.720 173.005 978.520 195.740 ;
        RECT 982.520 173.005 1030.720 195.740 ;
        RECT 754.520 45.435 1030.720 173.005 ;
        RECT 754.520 40.640 807.520 45.435 ;
        RECT 811.520 40.640 859.720 45.435 ;
        RECT 863.720 40.640 864.520 45.435 ;
        RECT 868.520 40.640 916.720 45.435 ;
        RECT 920.720 40.640 921.520 45.435 ;
        RECT 925.520 40.640 973.720 45.435 ;
        RECT 977.720 40.640 1030.720 45.435 ;
        RECT 1034.720 40.640 1035.520 2672.240 ;
        RECT 1039.520 2672.205 1092.520 2672.240 ;
        RECT 1096.520 2672.205 1144.720 2672.240 ;
        RECT 1148.720 2672.205 1149.520 2672.240 ;
        RECT 1153.520 2672.205 1201.720 2672.240 ;
        RECT 1205.720 2672.205 1206.520 2672.240 ;
        RECT 1210.520 2672.205 1258.720 2672.240 ;
        RECT 1262.720 2672.205 1315.720 2672.240 ;
        RECT 1039.520 2403.195 1315.720 2672.205 ;
        RECT 1039.520 2400.740 1092.520 2403.195 ;
        RECT 1039.520 2367.140 1087.720 2400.740 ;
        RECT 1091.720 2367.140 1092.520 2400.740 ;
        RECT 1039.520 2365.365 1092.520 2367.140 ;
        RECT 1096.520 2365.365 1144.720 2403.195 ;
        RECT 1148.720 2365.365 1149.520 2403.195 ;
        RECT 1153.520 2365.365 1201.720 2403.195 ;
        RECT 1205.720 2365.365 1206.520 2403.195 ;
        RECT 1210.520 2365.365 1258.720 2403.195 ;
        RECT 1262.720 2400.740 1315.720 2403.195 ;
        RECT 1262.720 2367.140 1263.520 2400.740 ;
        RECT 1267.520 2367.140 1315.720 2400.740 ;
        RECT 1262.720 2365.365 1315.720 2367.140 ;
        RECT 1039.520 2087.515 1315.720 2365.365 ;
        RECT 1039.520 2085.740 1092.520 2087.515 ;
        RECT 1039.520 2052.140 1087.720 2085.740 ;
        RECT 1091.720 2052.140 1092.520 2085.740 ;
        RECT 1039.520 2050.365 1092.520 2052.140 ;
        RECT 1096.520 2050.365 1144.720 2087.515 ;
        RECT 1148.720 2050.365 1149.520 2087.515 ;
        RECT 1153.520 2050.365 1201.720 2087.515 ;
        RECT 1205.720 2050.365 1206.520 2087.515 ;
        RECT 1210.520 2050.365 1258.720 2087.515 ;
        RECT 1262.720 2085.740 1315.720 2087.515 ;
        RECT 1262.720 2052.140 1263.520 2085.740 ;
        RECT 1267.520 2052.140 1315.720 2085.740 ;
        RECT 1262.720 2050.365 1315.720 2052.140 ;
        RECT 1039.520 1772.515 1315.720 2050.365 ;
        RECT 1039.520 1770.740 1092.520 1772.515 ;
        RECT 1039.520 1737.140 1087.720 1770.740 ;
        RECT 1091.720 1737.140 1092.520 1770.740 ;
        RECT 1039.520 1735.365 1092.520 1737.140 ;
        RECT 1096.520 1735.365 1144.720 1772.515 ;
        RECT 1148.720 1735.365 1149.520 1772.515 ;
        RECT 1153.520 1735.365 1201.720 1772.515 ;
        RECT 1205.720 1735.365 1206.520 1772.515 ;
        RECT 1210.520 1735.365 1258.720 1772.515 ;
        RECT 1262.720 1770.740 1315.720 1772.515 ;
        RECT 1262.720 1737.140 1263.520 1770.740 ;
        RECT 1267.520 1737.140 1315.720 1770.740 ;
        RECT 1262.720 1735.365 1315.720 1737.140 ;
        RECT 1039.520 1457.515 1315.720 1735.365 ;
        RECT 1039.520 1455.740 1092.520 1457.515 ;
        RECT 1039.520 1422.140 1087.720 1455.740 ;
        RECT 1091.720 1422.140 1092.520 1455.740 ;
        RECT 1039.520 1420.365 1092.520 1422.140 ;
        RECT 1096.520 1420.365 1144.720 1457.515 ;
        RECT 1148.720 1420.365 1149.520 1457.515 ;
        RECT 1153.520 1420.365 1201.720 1457.515 ;
        RECT 1205.720 1420.365 1206.520 1457.515 ;
        RECT 1210.520 1420.365 1258.720 1457.515 ;
        RECT 1262.720 1455.740 1315.720 1457.515 ;
        RECT 1262.720 1422.140 1263.520 1455.740 ;
        RECT 1267.520 1422.140 1315.720 1455.740 ;
        RECT 1262.720 1420.365 1315.720 1422.140 ;
        RECT 1039.520 1142.515 1315.720 1420.365 ;
        RECT 1039.520 1140.740 1092.520 1142.515 ;
        RECT 1039.520 1107.140 1087.720 1140.740 ;
        RECT 1091.720 1107.140 1092.520 1140.740 ;
        RECT 1039.520 1105.365 1092.520 1107.140 ;
        RECT 1096.520 1105.365 1144.720 1142.515 ;
        RECT 1148.720 1105.365 1149.520 1142.515 ;
        RECT 1153.520 1105.365 1201.720 1142.515 ;
        RECT 1205.720 1105.365 1206.520 1142.515 ;
        RECT 1210.520 1105.365 1258.720 1142.515 ;
        RECT 1262.720 1140.740 1315.720 1142.515 ;
        RECT 1262.720 1107.140 1263.520 1140.740 ;
        RECT 1267.520 1107.140 1315.720 1140.740 ;
        RECT 1262.720 1105.365 1315.720 1107.140 ;
        RECT 1039.520 827.515 1315.720 1105.365 ;
        RECT 1039.520 825.740 1092.520 827.515 ;
        RECT 1039.520 792.140 1087.720 825.740 ;
        RECT 1091.720 792.140 1092.520 825.740 ;
        RECT 1039.520 790.365 1092.520 792.140 ;
        RECT 1096.520 790.365 1144.720 827.515 ;
        RECT 1148.720 790.365 1149.520 827.515 ;
        RECT 1153.520 790.365 1201.720 827.515 ;
        RECT 1205.720 790.365 1206.520 827.515 ;
        RECT 1210.520 790.365 1258.720 827.515 ;
        RECT 1262.720 825.740 1315.720 827.515 ;
        RECT 1262.720 792.140 1263.520 825.740 ;
        RECT 1267.520 792.140 1315.720 825.740 ;
        RECT 1262.720 790.365 1315.720 792.140 ;
        RECT 1039.520 512.515 1315.720 790.365 ;
        RECT 1039.520 510.740 1092.520 512.515 ;
        RECT 1039.520 477.140 1087.720 510.740 ;
        RECT 1091.720 477.140 1092.520 510.740 ;
        RECT 1039.520 475.365 1092.520 477.140 ;
        RECT 1096.520 475.365 1144.720 512.515 ;
        RECT 1148.720 475.365 1149.520 512.515 ;
        RECT 1153.520 475.365 1201.720 512.515 ;
        RECT 1205.720 475.365 1206.520 512.515 ;
        RECT 1210.520 475.365 1258.720 512.515 ;
        RECT 1262.720 510.740 1315.720 512.515 ;
        RECT 1262.720 477.140 1263.520 510.740 ;
        RECT 1267.520 477.140 1315.720 510.740 ;
        RECT 1262.720 475.365 1315.720 477.140 ;
        RECT 1039.520 197.515 1315.720 475.365 ;
        RECT 1039.520 195.740 1092.520 197.515 ;
        RECT 1039.520 173.005 1087.720 195.740 ;
        RECT 1091.720 173.005 1092.520 195.740 ;
        RECT 1096.520 173.005 1144.720 197.515 ;
        RECT 1148.720 173.005 1149.520 197.515 ;
        RECT 1153.520 173.005 1201.720 197.515 ;
        RECT 1205.720 173.005 1206.520 197.515 ;
        RECT 1210.520 173.005 1258.720 197.515 ;
        RECT 1262.720 195.740 1315.720 197.515 ;
        RECT 1262.720 173.005 1263.520 195.740 ;
        RECT 1267.520 173.005 1315.720 195.740 ;
        RECT 1039.520 45.435 1315.720 173.005 ;
        RECT 1039.520 40.640 1092.520 45.435 ;
        RECT 1096.520 40.640 1144.720 45.435 ;
        RECT 1148.720 40.640 1149.520 45.435 ;
        RECT 1153.520 40.640 1201.720 45.435 ;
        RECT 1205.720 40.640 1206.520 45.435 ;
        RECT 1210.520 40.640 1258.720 45.435 ;
        RECT 1262.720 40.640 1315.720 45.435 ;
        RECT 1319.720 40.640 1320.520 2672.240 ;
        RECT 1324.520 2672.205 1377.520 2672.240 ;
        RECT 1381.520 2672.205 1429.720 2672.240 ;
        RECT 1433.720 2672.205 1434.520 2672.240 ;
        RECT 1438.520 2672.205 1486.720 2672.240 ;
        RECT 1490.720 2672.205 1491.520 2672.240 ;
        RECT 1495.520 2672.205 1543.720 2672.240 ;
        RECT 1547.720 2672.205 1600.720 2672.240 ;
        RECT 1324.520 2403.195 1600.720 2672.205 ;
        RECT 1324.520 2400.740 1377.520 2403.195 ;
        RECT 1324.520 2367.140 1372.720 2400.740 ;
        RECT 1376.720 2367.140 1377.520 2400.740 ;
        RECT 1324.520 2365.365 1377.520 2367.140 ;
        RECT 1381.520 2365.365 1429.720 2403.195 ;
        RECT 1433.720 2365.365 1434.520 2403.195 ;
        RECT 1438.520 2365.365 1486.720 2403.195 ;
        RECT 1490.720 2365.365 1491.520 2403.195 ;
        RECT 1495.520 2365.365 1543.720 2403.195 ;
        RECT 1547.720 2400.740 1600.720 2403.195 ;
        RECT 1547.720 2367.140 1548.520 2400.740 ;
        RECT 1552.520 2367.140 1600.720 2400.740 ;
        RECT 1547.720 2365.365 1600.720 2367.140 ;
        RECT 1324.520 2087.515 1600.720 2365.365 ;
        RECT 1324.520 2085.740 1377.520 2087.515 ;
        RECT 1324.520 2052.140 1372.720 2085.740 ;
        RECT 1376.720 2052.140 1377.520 2085.740 ;
        RECT 1324.520 2050.365 1377.520 2052.140 ;
        RECT 1381.520 2050.365 1429.720 2087.515 ;
        RECT 1433.720 2050.365 1434.520 2087.515 ;
        RECT 1438.520 2050.365 1486.720 2087.515 ;
        RECT 1490.720 2050.365 1491.520 2087.515 ;
        RECT 1495.520 2050.365 1543.720 2087.515 ;
        RECT 1547.720 2085.740 1600.720 2087.515 ;
        RECT 1547.720 2052.140 1548.520 2085.740 ;
        RECT 1552.520 2052.140 1600.720 2085.740 ;
        RECT 1547.720 2050.365 1600.720 2052.140 ;
        RECT 1324.520 1772.515 1600.720 2050.365 ;
        RECT 1324.520 1770.740 1377.520 1772.515 ;
        RECT 1324.520 1737.140 1372.720 1770.740 ;
        RECT 1376.720 1737.140 1377.520 1770.740 ;
        RECT 1324.520 1735.365 1377.520 1737.140 ;
        RECT 1381.520 1735.365 1429.720 1772.515 ;
        RECT 1433.720 1735.365 1434.520 1772.515 ;
        RECT 1438.520 1735.365 1486.720 1772.515 ;
        RECT 1490.720 1735.365 1491.520 1772.515 ;
        RECT 1495.520 1735.365 1543.720 1772.515 ;
        RECT 1547.720 1770.740 1600.720 1772.515 ;
        RECT 1547.720 1737.140 1548.520 1770.740 ;
        RECT 1552.520 1737.140 1600.720 1770.740 ;
        RECT 1547.720 1735.365 1600.720 1737.140 ;
        RECT 1324.520 1457.515 1600.720 1735.365 ;
        RECT 1324.520 1455.740 1377.520 1457.515 ;
        RECT 1324.520 1422.140 1372.720 1455.740 ;
        RECT 1376.720 1422.140 1377.520 1455.740 ;
        RECT 1324.520 1420.365 1377.520 1422.140 ;
        RECT 1381.520 1420.365 1429.720 1457.515 ;
        RECT 1433.720 1420.365 1434.520 1457.515 ;
        RECT 1438.520 1420.365 1486.720 1457.515 ;
        RECT 1490.720 1420.365 1491.520 1457.515 ;
        RECT 1495.520 1420.365 1543.720 1457.515 ;
        RECT 1547.720 1455.740 1600.720 1457.515 ;
        RECT 1547.720 1422.140 1548.520 1455.740 ;
        RECT 1552.520 1422.140 1600.720 1455.740 ;
        RECT 1547.720 1420.365 1600.720 1422.140 ;
        RECT 1324.520 1142.515 1600.720 1420.365 ;
        RECT 1324.520 1140.740 1377.520 1142.515 ;
        RECT 1324.520 1107.140 1372.720 1140.740 ;
        RECT 1376.720 1107.140 1377.520 1140.740 ;
        RECT 1324.520 1105.365 1377.520 1107.140 ;
        RECT 1381.520 1105.365 1429.720 1142.515 ;
        RECT 1433.720 1105.365 1434.520 1142.515 ;
        RECT 1438.520 1105.365 1486.720 1142.515 ;
        RECT 1490.720 1105.365 1491.520 1142.515 ;
        RECT 1495.520 1105.365 1543.720 1142.515 ;
        RECT 1547.720 1140.740 1600.720 1142.515 ;
        RECT 1547.720 1107.140 1548.520 1140.740 ;
        RECT 1552.520 1107.140 1600.720 1140.740 ;
        RECT 1547.720 1105.365 1600.720 1107.140 ;
        RECT 1324.520 827.515 1600.720 1105.365 ;
        RECT 1324.520 825.740 1377.520 827.515 ;
        RECT 1324.520 792.140 1372.720 825.740 ;
        RECT 1376.720 792.140 1377.520 825.740 ;
        RECT 1324.520 790.365 1377.520 792.140 ;
        RECT 1381.520 790.365 1429.720 827.515 ;
        RECT 1433.720 790.365 1434.520 827.515 ;
        RECT 1438.520 790.365 1486.720 827.515 ;
        RECT 1490.720 790.365 1491.520 827.515 ;
        RECT 1495.520 790.365 1543.720 827.515 ;
        RECT 1547.720 825.740 1600.720 827.515 ;
        RECT 1547.720 792.140 1548.520 825.740 ;
        RECT 1552.520 792.140 1600.720 825.740 ;
        RECT 1547.720 790.365 1600.720 792.140 ;
        RECT 1324.520 512.515 1600.720 790.365 ;
        RECT 1324.520 510.740 1377.520 512.515 ;
        RECT 1324.520 477.140 1372.720 510.740 ;
        RECT 1376.720 477.140 1377.520 510.740 ;
        RECT 1324.520 475.365 1377.520 477.140 ;
        RECT 1381.520 475.365 1429.720 512.515 ;
        RECT 1433.720 475.365 1434.520 512.515 ;
        RECT 1438.520 475.365 1486.720 512.515 ;
        RECT 1490.720 475.365 1491.520 512.515 ;
        RECT 1495.520 475.365 1543.720 512.515 ;
        RECT 1547.720 510.740 1600.720 512.515 ;
        RECT 1547.720 477.140 1548.520 510.740 ;
        RECT 1552.520 477.140 1600.720 510.740 ;
        RECT 1547.720 475.365 1600.720 477.140 ;
        RECT 1324.520 197.515 1600.720 475.365 ;
        RECT 1324.520 195.740 1377.520 197.515 ;
        RECT 1324.520 173.005 1372.720 195.740 ;
        RECT 1376.720 173.005 1377.520 195.740 ;
        RECT 1381.520 173.005 1429.720 197.515 ;
        RECT 1433.720 173.005 1434.520 197.515 ;
        RECT 1438.520 173.005 1486.720 197.515 ;
        RECT 1490.720 173.005 1491.520 197.515 ;
        RECT 1495.520 173.005 1543.720 197.515 ;
        RECT 1547.720 195.740 1600.720 197.515 ;
        RECT 1547.720 173.005 1548.520 195.740 ;
        RECT 1552.520 173.005 1600.720 195.740 ;
        RECT 1324.520 45.435 1600.720 173.005 ;
        RECT 1324.520 40.640 1377.520 45.435 ;
        RECT 1381.520 40.640 1429.720 45.435 ;
        RECT 1433.720 40.640 1434.520 45.435 ;
        RECT 1438.520 40.640 1486.720 45.435 ;
        RECT 1490.720 40.640 1491.520 45.435 ;
        RECT 1495.520 40.640 1543.720 45.435 ;
        RECT 1547.720 40.640 1600.720 45.435 ;
        RECT 1604.720 40.640 1605.520 2672.240 ;
        RECT 1609.520 2672.205 1662.520 2672.240 ;
        RECT 1666.520 2672.205 1714.720 2672.240 ;
        RECT 1718.720 2672.205 1719.520 2672.240 ;
        RECT 1723.520 2672.205 1771.720 2672.240 ;
        RECT 1775.720 2672.205 1776.520 2672.240 ;
        RECT 1780.520 2672.205 1828.720 2672.240 ;
        RECT 1832.720 2672.205 1885.720 2672.240 ;
        RECT 1609.520 2403.195 1885.720 2672.205 ;
        RECT 1609.520 2400.740 1662.520 2403.195 ;
        RECT 1609.520 2367.140 1657.720 2400.740 ;
        RECT 1661.720 2367.140 1662.520 2400.740 ;
        RECT 1609.520 2365.365 1662.520 2367.140 ;
        RECT 1666.520 2365.365 1714.720 2403.195 ;
        RECT 1718.720 2365.365 1719.520 2403.195 ;
        RECT 1723.520 2365.365 1771.720 2403.195 ;
        RECT 1775.720 2365.365 1776.520 2403.195 ;
        RECT 1780.520 2365.365 1828.720 2403.195 ;
        RECT 1832.720 2400.740 1885.720 2403.195 ;
        RECT 1832.720 2367.140 1833.520 2400.740 ;
        RECT 1837.520 2367.140 1885.720 2400.740 ;
        RECT 1832.720 2365.365 1885.720 2367.140 ;
        RECT 1609.520 2087.515 1885.720 2365.365 ;
        RECT 1609.520 2085.740 1662.520 2087.515 ;
        RECT 1609.520 2052.140 1657.720 2085.740 ;
        RECT 1661.720 2052.140 1662.520 2085.740 ;
        RECT 1609.520 2050.365 1662.520 2052.140 ;
        RECT 1666.520 2050.365 1714.720 2087.515 ;
        RECT 1718.720 2050.365 1719.520 2087.515 ;
        RECT 1723.520 2050.365 1771.720 2087.515 ;
        RECT 1775.720 2050.365 1776.520 2087.515 ;
        RECT 1780.520 2050.365 1828.720 2087.515 ;
        RECT 1832.720 2085.740 1885.720 2087.515 ;
        RECT 1832.720 2052.140 1833.520 2085.740 ;
        RECT 1837.520 2052.140 1885.720 2085.740 ;
        RECT 1832.720 2050.365 1885.720 2052.140 ;
        RECT 1609.520 1772.515 1885.720 2050.365 ;
        RECT 1609.520 1770.740 1662.520 1772.515 ;
        RECT 1609.520 1737.140 1657.720 1770.740 ;
        RECT 1661.720 1737.140 1662.520 1770.740 ;
        RECT 1609.520 1735.365 1662.520 1737.140 ;
        RECT 1666.520 1735.365 1714.720 1772.515 ;
        RECT 1718.720 1735.365 1719.520 1772.515 ;
        RECT 1723.520 1735.365 1771.720 1772.515 ;
        RECT 1775.720 1735.365 1776.520 1772.515 ;
        RECT 1780.520 1735.365 1828.720 1772.515 ;
        RECT 1832.720 1770.740 1885.720 1772.515 ;
        RECT 1832.720 1737.140 1833.520 1770.740 ;
        RECT 1837.520 1737.140 1885.720 1770.740 ;
        RECT 1832.720 1735.365 1885.720 1737.140 ;
        RECT 1609.520 1457.515 1885.720 1735.365 ;
        RECT 1609.520 1455.740 1662.520 1457.515 ;
        RECT 1609.520 1422.140 1657.720 1455.740 ;
        RECT 1661.720 1422.140 1662.520 1455.740 ;
        RECT 1609.520 1420.365 1662.520 1422.140 ;
        RECT 1666.520 1420.365 1714.720 1457.515 ;
        RECT 1718.720 1420.365 1719.520 1457.515 ;
        RECT 1723.520 1420.365 1771.720 1457.515 ;
        RECT 1775.720 1420.365 1776.520 1457.515 ;
        RECT 1780.520 1420.365 1828.720 1457.515 ;
        RECT 1832.720 1455.740 1885.720 1457.515 ;
        RECT 1832.720 1422.140 1833.520 1455.740 ;
        RECT 1837.520 1422.140 1885.720 1455.740 ;
        RECT 1832.720 1420.365 1885.720 1422.140 ;
        RECT 1609.520 1142.515 1885.720 1420.365 ;
        RECT 1609.520 1140.740 1662.520 1142.515 ;
        RECT 1609.520 1107.140 1657.720 1140.740 ;
        RECT 1661.720 1107.140 1662.520 1140.740 ;
        RECT 1609.520 1105.365 1662.520 1107.140 ;
        RECT 1666.520 1105.365 1714.720 1142.515 ;
        RECT 1718.720 1105.365 1719.520 1142.515 ;
        RECT 1723.520 1105.365 1771.720 1142.515 ;
        RECT 1775.720 1105.365 1776.520 1142.515 ;
        RECT 1780.520 1105.365 1828.720 1142.515 ;
        RECT 1832.720 1140.740 1885.720 1142.515 ;
        RECT 1832.720 1107.140 1833.520 1140.740 ;
        RECT 1837.520 1107.140 1885.720 1140.740 ;
        RECT 1832.720 1105.365 1885.720 1107.140 ;
        RECT 1609.520 827.515 1885.720 1105.365 ;
        RECT 1609.520 825.740 1662.520 827.515 ;
        RECT 1609.520 792.140 1657.720 825.740 ;
        RECT 1661.720 792.140 1662.520 825.740 ;
        RECT 1609.520 790.365 1662.520 792.140 ;
        RECT 1666.520 790.365 1714.720 827.515 ;
        RECT 1718.720 790.365 1719.520 827.515 ;
        RECT 1723.520 790.365 1771.720 827.515 ;
        RECT 1775.720 790.365 1776.520 827.515 ;
        RECT 1780.520 790.365 1828.720 827.515 ;
        RECT 1832.720 825.740 1885.720 827.515 ;
        RECT 1832.720 792.140 1833.520 825.740 ;
        RECT 1837.520 792.140 1885.720 825.740 ;
        RECT 1832.720 790.365 1885.720 792.140 ;
        RECT 1609.520 512.515 1885.720 790.365 ;
        RECT 1609.520 510.740 1662.520 512.515 ;
        RECT 1609.520 477.140 1657.720 510.740 ;
        RECT 1661.720 477.140 1662.520 510.740 ;
        RECT 1609.520 475.365 1662.520 477.140 ;
        RECT 1666.520 475.365 1714.720 512.515 ;
        RECT 1718.720 475.365 1719.520 512.515 ;
        RECT 1723.520 475.365 1771.720 512.515 ;
        RECT 1775.720 475.365 1776.520 512.515 ;
        RECT 1780.520 475.365 1828.720 512.515 ;
        RECT 1832.720 510.740 1885.720 512.515 ;
        RECT 1832.720 477.140 1833.520 510.740 ;
        RECT 1837.520 477.140 1885.720 510.740 ;
        RECT 1832.720 475.365 1885.720 477.140 ;
        RECT 1609.520 197.515 1885.720 475.365 ;
        RECT 1609.520 195.740 1662.520 197.515 ;
        RECT 1609.520 173.005 1657.720 195.740 ;
        RECT 1661.720 173.005 1662.520 195.740 ;
        RECT 1666.520 173.005 1714.720 197.515 ;
        RECT 1718.720 173.005 1719.520 197.515 ;
        RECT 1723.520 173.005 1771.720 197.515 ;
        RECT 1775.720 173.005 1776.520 197.515 ;
        RECT 1780.520 173.005 1828.720 197.515 ;
        RECT 1832.720 195.740 1885.720 197.515 ;
        RECT 1832.720 173.005 1833.520 195.740 ;
        RECT 1837.520 173.005 1885.720 195.740 ;
        RECT 1609.520 45.435 1885.720 173.005 ;
        RECT 1609.520 40.640 1662.520 45.435 ;
        RECT 1666.520 40.640 1714.720 45.435 ;
        RECT 1718.720 40.640 1719.520 45.435 ;
        RECT 1723.520 40.640 1771.720 45.435 ;
        RECT 1775.720 40.640 1776.520 45.435 ;
        RECT 1780.520 40.640 1828.720 45.435 ;
        RECT 1832.720 40.640 1885.720 45.435 ;
        RECT 1889.720 40.640 1890.520 2672.240 ;
        RECT 1894.520 2672.205 1947.520 2672.240 ;
        RECT 1951.520 2672.205 1999.720 2672.240 ;
        RECT 2003.720 2672.205 2004.520 2672.240 ;
        RECT 2008.520 2672.205 2056.720 2672.240 ;
        RECT 2060.720 2672.205 2061.520 2672.240 ;
        RECT 2065.520 2672.205 2113.720 2672.240 ;
        RECT 2117.720 2672.205 2170.720 2672.240 ;
        RECT 1894.520 2403.195 2170.720 2672.205 ;
        RECT 1894.520 2400.740 1947.520 2403.195 ;
        RECT 1894.520 2367.140 1942.720 2400.740 ;
        RECT 1946.720 2367.140 1947.520 2400.740 ;
        RECT 1894.520 2365.365 1947.520 2367.140 ;
        RECT 1951.520 2365.365 1999.720 2403.195 ;
        RECT 2003.720 2365.365 2004.520 2403.195 ;
        RECT 2008.520 2365.365 2056.720 2403.195 ;
        RECT 2060.720 2365.365 2061.520 2403.195 ;
        RECT 2065.520 2365.365 2113.720 2403.195 ;
        RECT 2117.720 2400.740 2170.720 2403.195 ;
        RECT 2117.720 2367.140 2118.520 2400.740 ;
        RECT 2122.520 2367.140 2170.720 2400.740 ;
        RECT 2117.720 2365.365 2170.720 2367.140 ;
        RECT 1894.520 2087.515 2170.720 2365.365 ;
        RECT 1894.520 2085.740 1947.520 2087.515 ;
        RECT 1894.520 2052.140 1942.720 2085.740 ;
        RECT 1946.720 2052.140 1947.520 2085.740 ;
        RECT 1894.520 2050.365 1947.520 2052.140 ;
        RECT 1951.520 2050.365 1999.720 2087.515 ;
        RECT 2003.720 2050.365 2004.520 2087.515 ;
        RECT 2008.520 2050.365 2056.720 2087.515 ;
        RECT 2060.720 2050.365 2061.520 2087.515 ;
        RECT 2065.520 2050.365 2113.720 2087.515 ;
        RECT 2117.720 2085.740 2170.720 2087.515 ;
        RECT 2117.720 2052.140 2118.520 2085.740 ;
        RECT 2122.520 2052.140 2170.720 2085.740 ;
        RECT 2117.720 2050.365 2170.720 2052.140 ;
        RECT 1894.520 1772.515 2170.720 2050.365 ;
        RECT 1894.520 1770.740 1947.520 1772.515 ;
        RECT 1894.520 1737.140 1942.720 1770.740 ;
        RECT 1946.720 1737.140 1947.520 1770.740 ;
        RECT 1894.520 1735.365 1947.520 1737.140 ;
        RECT 1951.520 1735.365 1999.720 1772.515 ;
        RECT 2003.720 1735.365 2004.520 1772.515 ;
        RECT 2008.520 1735.365 2056.720 1772.515 ;
        RECT 2060.720 1735.365 2061.520 1772.515 ;
        RECT 2065.520 1735.365 2113.720 1772.515 ;
        RECT 2117.720 1770.740 2170.720 1772.515 ;
        RECT 2117.720 1737.140 2118.520 1770.740 ;
        RECT 2122.520 1737.140 2170.720 1770.740 ;
        RECT 2117.720 1735.365 2170.720 1737.140 ;
        RECT 1894.520 1457.515 2170.720 1735.365 ;
        RECT 1894.520 1455.740 1947.520 1457.515 ;
        RECT 1894.520 1422.140 1942.720 1455.740 ;
        RECT 1946.720 1422.140 1947.520 1455.740 ;
        RECT 1894.520 1420.365 1947.520 1422.140 ;
        RECT 1951.520 1420.365 1999.720 1457.515 ;
        RECT 2003.720 1420.365 2004.520 1457.515 ;
        RECT 2008.520 1420.365 2056.720 1457.515 ;
        RECT 2060.720 1420.365 2061.520 1457.515 ;
        RECT 2065.520 1420.365 2113.720 1457.515 ;
        RECT 2117.720 1455.740 2170.720 1457.515 ;
        RECT 2117.720 1422.140 2118.520 1455.740 ;
        RECT 2122.520 1422.140 2170.720 1455.740 ;
        RECT 2117.720 1420.365 2170.720 1422.140 ;
        RECT 1894.520 1142.515 2170.720 1420.365 ;
        RECT 1894.520 1140.740 1947.520 1142.515 ;
        RECT 1894.520 1107.140 1942.720 1140.740 ;
        RECT 1946.720 1107.140 1947.520 1140.740 ;
        RECT 1894.520 1105.365 1947.520 1107.140 ;
        RECT 1951.520 1105.365 1999.720 1142.515 ;
        RECT 2003.720 1105.365 2004.520 1142.515 ;
        RECT 2008.520 1105.365 2056.720 1142.515 ;
        RECT 2060.720 1105.365 2061.520 1142.515 ;
        RECT 2065.520 1105.365 2113.720 1142.515 ;
        RECT 2117.720 1140.740 2170.720 1142.515 ;
        RECT 2117.720 1107.140 2118.520 1140.740 ;
        RECT 2122.520 1107.140 2170.720 1140.740 ;
        RECT 2117.720 1105.365 2170.720 1107.140 ;
        RECT 1894.520 827.515 2170.720 1105.365 ;
        RECT 1894.520 825.740 1947.520 827.515 ;
        RECT 1894.520 792.140 1942.720 825.740 ;
        RECT 1946.720 792.140 1947.520 825.740 ;
        RECT 1894.520 790.365 1947.520 792.140 ;
        RECT 1951.520 790.365 1999.720 827.515 ;
        RECT 2003.720 790.365 2004.520 827.515 ;
        RECT 2008.520 790.365 2056.720 827.515 ;
        RECT 2060.720 790.365 2061.520 827.515 ;
        RECT 2065.520 790.365 2113.720 827.515 ;
        RECT 2117.720 825.740 2170.720 827.515 ;
        RECT 2117.720 792.140 2118.520 825.740 ;
        RECT 2122.520 792.140 2170.720 825.740 ;
        RECT 2117.720 790.365 2170.720 792.140 ;
        RECT 1894.520 512.515 2170.720 790.365 ;
        RECT 1894.520 510.740 1947.520 512.515 ;
        RECT 1894.520 477.140 1942.720 510.740 ;
        RECT 1946.720 477.140 1947.520 510.740 ;
        RECT 1894.520 475.365 1947.520 477.140 ;
        RECT 1951.520 475.365 1999.720 512.515 ;
        RECT 2003.720 475.365 2004.520 512.515 ;
        RECT 2008.520 475.365 2056.720 512.515 ;
        RECT 2060.720 475.365 2061.520 512.515 ;
        RECT 2065.520 475.365 2113.720 512.515 ;
        RECT 2117.720 510.740 2170.720 512.515 ;
        RECT 2117.720 477.140 2118.520 510.740 ;
        RECT 2122.520 477.140 2170.720 510.740 ;
        RECT 2117.720 475.365 2170.720 477.140 ;
        RECT 1894.520 197.515 2170.720 475.365 ;
        RECT 1894.520 195.740 1947.520 197.515 ;
        RECT 1894.520 173.005 1942.720 195.740 ;
        RECT 1946.720 173.005 1947.520 195.740 ;
        RECT 1951.520 173.005 1999.720 197.515 ;
        RECT 2003.720 173.005 2004.520 197.515 ;
        RECT 2008.520 173.005 2056.720 197.515 ;
        RECT 2060.720 173.005 2061.520 197.515 ;
        RECT 2065.520 173.005 2113.720 197.515 ;
        RECT 2117.720 195.740 2170.720 197.515 ;
        RECT 2117.720 173.005 2118.520 195.740 ;
        RECT 2122.520 173.005 2170.720 195.740 ;
        RECT 1894.520 45.435 2170.720 173.005 ;
        RECT 1894.520 40.640 1947.520 45.435 ;
        RECT 1951.520 40.640 1999.720 45.435 ;
        RECT 2003.720 40.640 2004.520 45.435 ;
        RECT 2008.520 40.640 2056.720 45.435 ;
        RECT 2060.720 40.640 2061.520 45.435 ;
        RECT 2065.520 40.640 2113.720 45.435 ;
        RECT 2117.720 40.640 2170.720 45.435 ;
        RECT 2174.720 40.640 2175.520 2672.240 ;
        RECT 2179.520 2655.885 2232.520 2672.240 ;
        RECT 2236.520 2655.885 2284.720 2672.240 ;
        RECT 2288.720 2655.885 2289.520 2672.240 ;
        RECT 2293.520 2655.885 2341.720 2672.240 ;
        RECT 2345.720 2655.885 2346.520 2672.240 ;
        RECT 2350.520 2655.885 2398.720 2672.240 ;
        RECT 2402.720 2655.885 2431.320 2672.240 ;
        RECT 2179.520 2402.515 2431.320 2655.885 ;
        RECT 2179.520 2400.740 2232.520 2402.515 ;
        RECT 2179.520 2367.140 2227.720 2400.740 ;
        RECT 2231.720 2367.140 2232.520 2400.740 ;
        RECT 2179.520 2365.365 2232.520 2367.140 ;
        RECT 2236.520 2365.365 2284.720 2402.515 ;
        RECT 2288.720 2365.365 2289.520 2402.515 ;
        RECT 2293.520 2365.365 2341.720 2402.515 ;
        RECT 2345.720 2365.365 2346.520 2402.515 ;
        RECT 2350.520 2365.365 2398.720 2402.515 ;
        RECT 2402.720 2400.740 2431.320 2402.515 ;
        RECT 2402.720 2367.140 2403.520 2400.740 ;
        RECT 2407.520 2367.140 2431.320 2400.740 ;
        RECT 2402.720 2365.365 2431.320 2367.140 ;
        RECT 2179.520 2087.515 2431.320 2365.365 ;
        RECT 2179.520 2085.740 2232.520 2087.515 ;
        RECT 2179.520 2052.140 2227.720 2085.740 ;
        RECT 2231.720 2052.140 2232.520 2085.740 ;
        RECT 2179.520 2050.365 2232.520 2052.140 ;
        RECT 2236.520 2050.365 2284.720 2087.515 ;
        RECT 2288.720 2050.365 2289.520 2087.515 ;
        RECT 2293.520 2050.365 2341.720 2087.515 ;
        RECT 2345.720 2050.365 2346.520 2087.515 ;
        RECT 2350.520 2050.365 2398.720 2087.515 ;
        RECT 2402.720 2085.740 2431.320 2087.515 ;
        RECT 2402.720 2052.140 2403.520 2085.740 ;
        RECT 2407.520 2052.140 2431.320 2085.740 ;
        RECT 2402.720 2050.365 2431.320 2052.140 ;
        RECT 2179.520 1772.515 2431.320 2050.365 ;
        RECT 2179.520 1770.740 2232.520 1772.515 ;
        RECT 2179.520 1737.140 2227.720 1770.740 ;
        RECT 2231.720 1737.140 2232.520 1770.740 ;
        RECT 2179.520 1735.365 2232.520 1737.140 ;
        RECT 2236.520 1735.365 2284.720 1772.515 ;
        RECT 2288.720 1735.365 2289.520 1772.515 ;
        RECT 2293.520 1735.365 2341.720 1772.515 ;
        RECT 2345.720 1735.365 2346.520 1772.515 ;
        RECT 2350.520 1735.365 2398.720 1772.515 ;
        RECT 2402.720 1770.740 2431.320 1772.515 ;
        RECT 2402.720 1737.140 2403.520 1770.740 ;
        RECT 2407.520 1737.140 2431.320 1770.740 ;
        RECT 2402.720 1735.365 2431.320 1737.140 ;
        RECT 2179.520 1457.515 2431.320 1735.365 ;
        RECT 2179.520 1455.740 2232.520 1457.515 ;
        RECT 2179.520 1422.140 2227.720 1455.740 ;
        RECT 2231.720 1422.140 2232.520 1455.740 ;
        RECT 2179.520 1420.365 2232.520 1422.140 ;
        RECT 2236.520 1420.365 2284.720 1457.515 ;
        RECT 2288.720 1420.365 2289.520 1457.515 ;
        RECT 2293.520 1420.365 2341.720 1457.515 ;
        RECT 2345.720 1420.365 2346.520 1457.515 ;
        RECT 2350.520 1420.365 2398.720 1457.515 ;
        RECT 2402.720 1455.740 2431.320 1457.515 ;
        RECT 2402.720 1422.140 2403.520 1455.740 ;
        RECT 2407.520 1422.140 2431.320 1455.740 ;
        RECT 2402.720 1420.365 2431.320 1422.140 ;
        RECT 2179.520 1142.515 2431.320 1420.365 ;
        RECT 2179.520 1140.740 2232.520 1142.515 ;
        RECT 2179.520 1107.140 2227.720 1140.740 ;
        RECT 2231.720 1107.140 2232.520 1140.740 ;
        RECT 2179.520 1105.365 2232.520 1107.140 ;
        RECT 2236.520 1105.365 2284.720 1142.515 ;
        RECT 2288.720 1105.365 2289.520 1142.515 ;
        RECT 2293.520 1105.365 2341.720 1142.515 ;
        RECT 2345.720 1105.365 2346.520 1142.515 ;
        RECT 2350.520 1105.365 2398.720 1142.515 ;
        RECT 2402.720 1140.740 2431.320 1142.515 ;
        RECT 2402.720 1107.140 2403.520 1140.740 ;
        RECT 2407.520 1107.140 2431.320 1140.740 ;
        RECT 2402.720 1105.365 2431.320 1107.140 ;
        RECT 2179.520 827.515 2431.320 1105.365 ;
        RECT 2179.520 825.740 2232.520 827.515 ;
        RECT 2179.520 792.140 2227.720 825.740 ;
        RECT 2231.720 792.140 2232.520 825.740 ;
        RECT 2179.520 790.365 2232.520 792.140 ;
        RECT 2236.520 790.365 2284.720 827.515 ;
        RECT 2288.720 790.365 2289.520 827.515 ;
        RECT 2293.520 790.365 2341.720 827.515 ;
        RECT 2345.720 790.365 2346.520 827.515 ;
        RECT 2350.520 790.365 2398.720 827.515 ;
        RECT 2402.720 825.740 2431.320 827.515 ;
        RECT 2402.720 792.140 2403.520 825.740 ;
        RECT 2407.520 792.140 2431.320 825.740 ;
        RECT 2402.720 790.365 2431.320 792.140 ;
        RECT 2179.520 512.515 2431.320 790.365 ;
        RECT 2179.520 510.740 2232.520 512.515 ;
        RECT 2179.520 477.140 2227.720 510.740 ;
        RECT 2231.720 477.140 2232.520 510.740 ;
        RECT 2179.520 475.365 2232.520 477.140 ;
        RECT 2236.520 475.365 2284.720 512.515 ;
        RECT 2288.720 475.365 2289.520 512.515 ;
        RECT 2293.520 475.365 2341.720 512.515 ;
        RECT 2345.720 475.365 2346.520 512.515 ;
        RECT 2350.520 475.365 2398.720 512.515 ;
        RECT 2402.720 510.740 2431.320 512.515 ;
        RECT 2402.720 477.140 2403.520 510.740 ;
        RECT 2407.520 477.140 2431.320 510.740 ;
        RECT 2402.720 475.365 2431.320 477.140 ;
        RECT 2179.520 197.515 2431.320 475.365 ;
        RECT 2179.520 195.740 2232.520 197.515 ;
        RECT 2179.520 171.645 2227.720 195.740 ;
        RECT 2231.720 171.645 2232.520 195.740 ;
        RECT 2236.520 171.645 2284.720 197.515 ;
        RECT 2288.720 171.645 2289.520 197.515 ;
        RECT 2293.520 171.645 2341.720 197.515 ;
        RECT 2345.720 171.645 2346.520 197.515 ;
        RECT 2350.520 171.645 2398.720 197.515 ;
        RECT 2179.520 48.155 2398.720 171.645 ;
        RECT 2179.520 40.640 2232.520 48.155 ;
        RECT 2236.520 40.640 2284.720 48.155 ;
        RECT 2288.720 40.640 2289.520 48.155 ;
        RECT 2293.520 40.640 2341.720 48.155 ;
        RECT 2345.720 40.640 2346.520 48.155 ;
        RECT 2350.520 40.640 2398.720 48.155 ;
        RECT 2402.720 195.740 2431.320 197.515 ;
        RECT 2402.720 162.540 2403.520 195.740 ;
        RECT 2407.520 162.540 2431.320 195.740 ;
        RECT 2402.720 40.640 2431.320 162.540 ;
  END
END fpga_core
END LIBRARY

