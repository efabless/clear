magic
tech sky130A
magscale 1 2
timestamp 1656945640
<< viali >>
rect 9689 20553 9723 20587
rect 20361 20553 20395 20587
rect 20821 20553 20855 20587
rect 9873 20417 9907 20451
rect 16957 20417 16991 20451
rect 20637 20417 20671 20451
rect 17141 20213 17175 20247
rect 18797 20213 18831 20247
rect 19901 20213 19935 20247
rect 21189 20213 21223 20247
rect 5733 20009 5767 20043
rect 11713 20009 11747 20043
rect 18061 20009 18095 20043
rect 19349 20009 19383 20043
rect 7389 19941 7423 19975
rect 14841 19941 14875 19975
rect 17509 19941 17543 19975
rect 18521 19941 18555 19975
rect 19901 19941 19935 19975
rect 9229 19873 9263 19907
rect 10425 19873 10459 19907
rect 21005 19873 21039 19907
rect 4169 19805 4203 19839
rect 4721 19805 4755 19839
rect 5917 19805 5951 19839
rect 7205 19805 7239 19839
rect 9413 19805 9447 19839
rect 11529 19805 11563 19839
rect 14657 19805 14691 19839
rect 15209 19805 15243 19839
rect 16773 19805 16807 19839
rect 17325 19805 17359 19839
rect 17877 19805 17911 19839
rect 18705 19805 18739 19839
rect 19533 19805 19567 19839
rect 20085 19805 20119 19839
rect 21189 19805 21223 19839
rect 4997 19737 5031 19771
rect 10149 19737 10183 19771
rect 10793 19737 10827 19771
rect 4353 19669 4387 19703
rect 9781 19669 9815 19703
rect 10241 19669 10275 19703
rect 15393 19669 15427 19703
rect 16957 19669 16991 19703
rect 3893 19465 3927 19499
rect 9873 19465 9907 19499
rect 20729 19465 20763 19499
rect 7297 19397 7331 19431
rect 10701 19397 10735 19431
rect 12664 19397 12698 19431
rect 4077 19329 4111 19363
rect 7573 19329 7607 19363
rect 10057 19329 10091 19363
rect 10425 19329 10459 19363
rect 17325 19329 17359 19363
rect 17581 19329 17615 19363
rect 20913 19329 20947 19363
rect 12909 19261 12943 19295
rect 19717 19193 19751 19227
rect 11529 19125 11563 19159
rect 13277 19125 13311 19159
rect 18705 19125 18739 19159
rect 19073 19125 19107 19159
rect 20269 19125 20303 19159
rect 21281 19125 21315 19159
rect 16313 18921 16347 18955
rect 4077 18785 4111 18819
rect 8493 18785 8527 18819
rect 9137 18785 9171 18819
rect 2421 18717 2455 18751
rect 4261 18717 4295 18751
rect 5181 18717 5215 18751
rect 8309 18717 8343 18751
rect 8953 18717 8987 18751
rect 12081 18717 12115 18751
rect 12357 18717 12391 18751
rect 14197 18717 14231 18751
rect 14933 18717 14967 18751
rect 16681 18717 16715 18751
rect 18705 18717 18739 18751
rect 19349 18717 19383 18751
rect 19901 18717 19935 18751
rect 2145 18649 2179 18683
rect 4905 18649 4939 18683
rect 11814 18649 11848 18683
rect 12624 18649 12658 18683
rect 15200 18649 15234 18683
rect 18438 18649 18472 18683
rect 20146 18649 20180 18683
rect 7849 18581 7883 18615
rect 8217 18581 8251 18615
rect 9689 18581 9723 18615
rect 10701 18581 10735 18615
rect 13737 18581 13771 18615
rect 17325 18581 17359 18615
rect 21281 18581 21315 18615
rect 8677 18377 8711 18411
rect 9045 18377 9079 18411
rect 12081 18377 12115 18411
rect 14013 18377 14047 18411
rect 20637 18377 20671 18411
rect 4537 18309 4571 18343
rect 4813 18241 4847 18275
rect 6929 18241 6963 18275
rect 7573 18241 7607 18275
rect 9413 18241 9447 18275
rect 10057 18241 10091 18275
rect 13470 18241 13504 18275
rect 13737 18241 13771 18275
rect 18317 18241 18351 18275
rect 20269 18241 20303 18275
rect 20821 18241 20855 18275
rect 6653 18173 6687 18207
rect 6837 18173 6871 18207
rect 9505 18173 9539 18207
rect 9597 18173 9631 18207
rect 18061 18173 18095 18207
rect 19809 18105 19843 18139
rect 7297 18037 7331 18071
rect 12357 18037 12391 18071
rect 19441 18037 19475 18071
rect 21281 18037 21315 18071
rect 4537 17833 4571 17867
rect 9781 17833 9815 17867
rect 13185 17833 13219 17867
rect 13553 17833 13587 17867
rect 17233 17833 17267 17867
rect 6469 17765 6503 17799
rect 3893 17697 3927 17731
rect 5457 17697 5491 17731
rect 5641 17697 5675 17731
rect 9229 17697 9263 17731
rect 9321 17697 9355 17731
rect 10425 17697 10459 17731
rect 16865 17697 16899 17731
rect 11805 17629 11839 17663
rect 16609 17629 16643 17663
rect 20922 17629 20956 17663
rect 21189 17629 21223 17663
rect 4077 17561 4111 17595
rect 5365 17561 5399 17595
rect 6101 17561 6135 17595
rect 9413 17561 9447 17595
rect 10057 17561 10091 17595
rect 12050 17561 12084 17595
rect 4169 17493 4203 17527
rect 4997 17493 5031 17527
rect 15485 17493 15519 17527
rect 19809 17493 19843 17527
rect 4353 17289 4387 17323
rect 5273 17289 5307 17323
rect 10241 17289 10275 17323
rect 18337 17289 18371 17323
rect 5733 17221 5767 17255
rect 15761 17221 15795 17255
rect 5641 17153 5675 17187
rect 6377 17153 6411 17187
rect 6929 17153 6963 17187
rect 9873 17153 9907 17187
rect 10517 17153 10551 17187
rect 11529 17153 11563 17187
rect 11796 17153 11830 17187
rect 14372 17153 14406 17187
rect 17805 17153 17839 17187
rect 18061 17153 18095 17187
rect 20646 17153 20680 17187
rect 5917 17085 5951 17119
rect 9597 17085 9631 17119
rect 9781 17085 9815 17119
rect 13277 17085 13311 17119
rect 14105 17085 14139 17119
rect 20913 17085 20947 17119
rect 16681 17017 16715 17051
rect 19533 17017 19567 17051
rect 12909 16949 12943 16983
rect 15485 16949 15519 16983
rect 21281 16949 21315 16983
rect 6561 16745 6595 16779
rect 20913 16745 20947 16779
rect 4537 16609 4571 16643
rect 4721 16609 4755 16643
rect 6009 16609 6043 16643
rect 7297 16609 7331 16643
rect 7481 16609 7515 16643
rect 10241 16609 10275 16643
rect 11621 16609 11655 16643
rect 17693 16609 17727 16643
rect 21281 16609 21315 16643
rect 15218 16541 15252 16575
rect 15485 16541 15519 16575
rect 15853 16541 15887 16575
rect 18245 16541 18279 16575
rect 18521 16541 18555 16575
rect 20729 16541 20763 16575
rect 6193 16473 6227 16507
rect 9965 16473 9999 16507
rect 10609 16473 10643 16507
rect 11866 16473 11900 16507
rect 17426 16473 17460 16507
rect 4077 16405 4111 16439
rect 4445 16405 4479 16439
rect 5089 16405 5123 16439
rect 6101 16405 6135 16439
rect 6837 16405 6871 16439
rect 7205 16405 7239 16439
rect 7849 16405 7883 16439
rect 9597 16405 9631 16439
rect 10057 16405 10091 16439
rect 13001 16405 13035 16439
rect 13369 16405 13403 16439
rect 14105 16405 14139 16439
rect 16313 16405 16347 16439
rect 5641 16201 5675 16235
rect 8217 16201 8251 16235
rect 11897 16201 11931 16235
rect 17877 16201 17911 16235
rect 6653 16133 6687 16167
rect 7205 16065 7239 16099
rect 7757 16065 7791 16099
rect 7849 16065 7883 16099
rect 13010 16065 13044 16099
rect 21106 16065 21140 16099
rect 21373 16065 21407 16099
rect 7665 15997 7699 16031
rect 13277 15997 13311 16031
rect 8493 15861 8527 15895
rect 13553 15861 13587 15895
rect 19993 15861 20027 15895
rect 19349 15657 19383 15691
rect 21281 15657 21315 15691
rect 13021 15453 13055 15487
rect 13277 15453 13311 15487
rect 15669 15453 15703 15487
rect 18889 15453 18923 15487
rect 15914 15385 15948 15419
rect 18644 15385 18678 15419
rect 11897 15317 11931 15351
rect 13553 15317 13587 15351
rect 17049 15317 17083 15351
rect 17509 15317 17543 15351
rect 5273 15113 5307 15147
rect 5733 15113 5767 15147
rect 7021 15113 7055 15147
rect 8033 15113 8067 15147
rect 16773 15113 16807 15147
rect 17233 15113 17267 15147
rect 9505 15045 9539 15079
rect 15976 15045 16010 15079
rect 20922 15045 20956 15079
rect 5641 14977 5675 15011
rect 6929 14977 6963 15011
rect 16221 14977 16255 15011
rect 21189 14977 21223 15011
rect 5917 14909 5951 14943
rect 7205 14909 7239 14943
rect 6561 14773 6595 14807
rect 7665 14773 7699 14807
rect 14841 14773 14875 14807
rect 19809 14773 19843 14807
rect 11621 14569 11655 14603
rect 15853 14569 15887 14603
rect 21097 14569 21131 14603
rect 17509 14501 17543 14535
rect 5733 14433 5767 14467
rect 8033 14433 8067 14467
rect 9781 14433 9815 14467
rect 15485 14433 15519 14467
rect 18889 14433 18923 14467
rect 19349 14433 19383 14467
rect 9965 14365 9999 14399
rect 10057 14365 10091 14399
rect 10701 14365 10735 14399
rect 13001 14365 13035 14399
rect 19605 14365 19639 14399
rect 8217 14297 8251 14331
rect 8953 14297 8987 14331
rect 12756 14297 12790 14331
rect 15218 14297 15252 14331
rect 17233 14297 17267 14331
rect 18622 14297 18656 14331
rect 8125 14229 8159 14263
rect 8585 14229 8619 14263
rect 10425 14229 10459 14263
rect 13369 14229 13403 14263
rect 14105 14229 14139 14263
rect 20729 14229 20763 14263
rect 8217 14025 8251 14059
rect 9137 14025 9171 14059
rect 9597 14025 9631 14059
rect 10517 14025 10551 14059
rect 13553 14025 13587 14059
rect 19073 14025 19107 14059
rect 20821 14025 20855 14059
rect 7849 13957 7883 13991
rect 8585 13957 8619 13991
rect 9505 13957 9539 13991
rect 7205 13889 7239 13923
rect 7757 13889 7791 13923
rect 12173 13889 12207 13923
rect 12429 13889 12463 13923
rect 7665 13821 7699 13855
rect 9689 13821 9723 13855
rect 10149 13821 10183 13855
rect 13921 13821 13955 13855
rect 21281 13685 21315 13719
rect 5917 13481 5951 13515
rect 7389 13481 7423 13515
rect 9689 13481 9723 13515
rect 10885 13481 10919 13515
rect 13461 13481 13495 13515
rect 16405 13481 16439 13515
rect 21005 13481 21039 13515
rect 6469 13345 6503 13379
rect 9137 13345 9171 13379
rect 16129 13345 16163 13379
rect 20637 13345 20671 13379
rect 6561 13277 6595 13311
rect 6653 13277 6687 13311
rect 9229 13277 9263 13311
rect 11713 13277 11747 13311
rect 17978 13277 18012 13311
rect 18245 13277 18279 13311
rect 18613 13277 18647 13311
rect 21189 13277 21223 13311
rect 9321 13209 9355 13243
rect 9965 13209 9999 13243
rect 11980 13209 12014 13243
rect 15862 13209 15896 13243
rect 20370 13209 20404 13243
rect 7021 13141 7055 13175
rect 10425 13141 10459 13175
rect 13093 13141 13127 13175
rect 14749 13141 14783 13175
rect 16865 13141 16899 13175
rect 19257 13141 19291 13175
rect 10057 12937 10091 12971
rect 10425 12937 10459 12971
rect 10517 12937 10551 12971
rect 13461 12937 13495 12971
rect 18429 12937 18463 12971
rect 12826 12869 12860 12903
rect 13093 12801 13127 12835
rect 16681 12801 16715 12835
rect 16937 12801 16971 12835
rect 21106 12801 21140 12835
rect 21373 12801 21407 12835
rect 10701 12733 10735 12767
rect 19625 12665 19659 12699
rect 11713 12597 11747 12631
rect 18061 12597 18095 12631
rect 19073 12597 19107 12631
rect 19993 12597 20027 12631
rect 10057 12257 10091 12291
rect 10241 12189 10275 12223
rect 21281 12189 21315 12223
rect 21014 12121 21048 12155
rect 6009 12053 6043 12087
rect 19533 12053 19567 12087
rect 19901 12053 19935 12087
rect 6745 11849 6779 11883
rect 7113 11849 7147 11883
rect 18981 11849 19015 11883
rect 6653 11781 6687 11815
rect 14125 11713 14159 11747
rect 14381 11713 14415 11747
rect 18438 11713 18472 11747
rect 20094 11713 20128 11747
rect 20361 11713 20395 11747
rect 20637 11713 20671 11747
rect 21281 11713 21315 11747
rect 6561 11645 6595 11679
rect 18705 11645 18739 11679
rect 13001 11509 13035 11543
rect 14749 11509 14783 11543
rect 17325 11509 17359 11543
rect 7389 11305 7423 11339
rect 10149 11305 10183 11339
rect 15945 11305 15979 11339
rect 20637 11305 20671 11339
rect 20913 11305 20947 11339
rect 15485 11237 15519 11271
rect 9597 11169 9631 11203
rect 9689 11101 9723 11135
rect 12725 11101 12759 11135
rect 13093 11101 13127 11135
rect 14105 11101 14139 11135
rect 17058 11101 17092 11135
rect 17325 11101 17359 11135
rect 17601 11101 17635 11135
rect 18797 11101 18831 11135
rect 19257 11101 19291 11135
rect 19513 11101 19547 11135
rect 9781 11033 9815 11067
rect 10425 11033 10459 11067
rect 12458 11033 12492 11067
rect 14350 11033 14384 11067
rect 11345 10965 11379 10999
rect 6837 10761 6871 10795
rect 7573 10761 7607 10795
rect 7941 10761 7975 10795
rect 13277 10761 13311 10795
rect 15669 10761 15703 10795
rect 15945 10761 15979 10795
rect 19809 10761 19843 10795
rect 8033 10693 8067 10727
rect 18521 10693 18555 10727
rect 6929 10625 6963 10659
rect 11529 10625 11563 10659
rect 11785 10625 11819 10659
rect 14758 10625 14792 10659
rect 15025 10625 15059 10659
rect 17978 10625 18012 10659
rect 18245 10625 18279 10659
rect 20922 10625 20956 10659
rect 21189 10625 21223 10659
rect 6745 10557 6779 10591
rect 8217 10557 8251 10591
rect 9321 10557 9355 10591
rect 12909 10489 12943 10523
rect 7297 10421 7331 10455
rect 8585 10421 8619 10455
rect 13645 10421 13679 10455
rect 16865 10421 16899 10455
rect 13277 10217 13311 10251
rect 15209 10217 15243 10251
rect 21281 10217 21315 10251
rect 7113 10081 7147 10115
rect 9229 10081 9263 10115
rect 10425 10081 10459 10115
rect 13001 10081 13035 10115
rect 16589 10081 16623 10115
rect 17233 10081 17267 10115
rect 8125 10013 8159 10047
rect 9413 10013 9447 10047
rect 10149 10013 10183 10047
rect 12745 10013 12779 10047
rect 16333 10013 16367 10047
rect 8401 9945 8435 9979
rect 9321 9877 9355 9911
rect 9781 9877 9815 9911
rect 11621 9877 11655 9911
rect 16865 9877 16899 9911
rect 7389 9605 7423 9639
rect 8217 9605 8251 9639
rect 8125 9537 8159 9571
rect 8769 9537 8803 9571
rect 12265 9537 12299 9571
rect 15209 9537 15243 9571
rect 15485 9537 15519 9571
rect 19717 9537 19751 9571
rect 20545 9537 20579 9571
rect 21373 9537 21407 9571
rect 8401 9469 8435 9503
rect 15025 9469 15059 9503
rect 7757 9401 7791 9435
rect 12449 9401 12483 9435
rect 15669 9401 15703 9435
rect 19901 9401 19935 9435
rect 20729 9401 20763 9435
rect 21189 9333 21223 9367
rect 7021 9129 7055 9163
rect 14197 9129 14231 9163
rect 15301 9129 15335 9163
rect 17233 9129 17267 9163
rect 19441 9129 19475 9163
rect 20453 9129 20487 9163
rect 6193 9061 6227 9095
rect 5549 8993 5583 9027
rect 5733 8993 5767 9027
rect 9229 8993 9263 9027
rect 13093 8993 13127 9027
rect 15945 8993 15979 9027
rect 17877 8993 17911 9027
rect 8953 8925 8987 8959
rect 13369 8925 13403 8959
rect 14565 8925 14599 8959
rect 15761 8925 15795 8959
rect 16865 8925 16899 8959
rect 17693 8925 17727 8959
rect 19257 8925 19291 8959
rect 19809 8925 19843 8959
rect 20637 8925 20671 8959
rect 21373 8925 21407 8959
rect 5825 8857 5859 8891
rect 6469 8857 6503 8891
rect 14841 8857 14875 8891
rect 12449 8789 12483 8823
rect 15669 8789 15703 8823
rect 16405 8789 16439 8823
rect 17601 8789 17635 8823
rect 18337 8789 18371 8823
rect 19993 8789 20027 8823
rect 21005 8789 21039 8823
rect 6745 8585 6779 8619
rect 7389 8585 7423 8619
rect 9229 8585 9263 8619
rect 9873 8585 9907 8619
rect 11805 8585 11839 8619
rect 12265 8585 12299 8619
rect 13277 8585 13311 8619
rect 15117 8585 15151 8619
rect 17509 8585 17543 8619
rect 18061 8585 18095 8619
rect 19257 8585 19291 8619
rect 19901 8585 19935 8619
rect 20453 8585 20487 8619
rect 10333 8517 10367 8551
rect 14749 8517 14783 8551
rect 15669 8517 15703 8551
rect 7481 8449 7515 8483
rect 10241 8449 10275 8483
rect 10885 8449 10919 8483
rect 11897 8449 11931 8483
rect 12909 8449 12943 8483
rect 13553 8449 13587 8483
rect 15945 8449 15979 8483
rect 17417 8449 17451 8483
rect 18429 8449 18463 8483
rect 19073 8449 19107 8483
rect 20085 8449 20119 8483
rect 20637 8449 20671 8483
rect 7297 8381 7331 8415
rect 8953 8381 8987 8415
rect 9137 8381 9171 8415
rect 10425 8381 10459 8415
rect 11621 8381 11655 8415
rect 12725 8381 12759 8415
rect 12817 8381 12851 8415
rect 14473 8381 14507 8415
rect 14657 8381 14691 8415
rect 17693 8381 17727 8415
rect 18521 8381 18555 8415
rect 18705 8381 18739 8415
rect 8125 8313 8159 8347
rect 17049 8313 17083 8347
rect 21005 8313 21039 8347
rect 21373 8313 21407 8347
rect 7849 8245 7883 8279
rect 9597 8245 9631 8279
rect 8309 8041 8343 8075
rect 10701 8041 10735 8075
rect 17049 8041 17083 8075
rect 19349 8041 19383 8075
rect 16773 7973 16807 8007
rect 18521 7973 18555 8007
rect 7665 7905 7699 7939
rect 7849 7905 7883 7939
rect 12173 7905 12207 7939
rect 17509 7905 17543 7939
rect 17693 7905 17727 7939
rect 18061 7905 18095 7939
rect 9413 7837 9447 7871
rect 9689 7837 9723 7871
rect 20913 7837 20947 7871
rect 17417 7769 17451 7803
rect 7941 7701 7975 7735
rect 20729 7701 20763 7735
rect 21281 7701 21315 7735
rect 7757 7497 7791 7531
rect 8217 7497 8251 7531
rect 14657 7497 14691 7531
rect 20177 7497 20211 7531
rect 7849 7429 7883 7463
rect 8861 7429 8895 7463
rect 19349 7429 19383 7463
rect 8493 7361 8527 7395
rect 10517 7361 10551 7395
rect 14473 7361 14507 7395
rect 19073 7361 19107 7395
rect 19993 7361 20027 7395
rect 21097 7361 21131 7395
rect 7573 7293 7607 7327
rect 10333 7293 10367 7327
rect 11529 7293 11563 7327
rect 17969 7293 18003 7327
rect 20913 7225 20947 7259
rect 7481 6817 7515 6851
rect 8033 6817 8067 6851
rect 9137 6817 9171 6851
rect 11437 6817 11471 6851
rect 15209 6817 15243 6851
rect 8125 6749 8159 6783
rect 10057 6749 10091 6783
rect 11253 6749 11287 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 19257 6749 19291 6783
rect 20085 6749 20119 6783
rect 21097 6749 21131 6783
rect 8217 6613 8251 6647
rect 8585 6613 8619 6647
rect 9229 6613 9263 6647
rect 9321 6613 9355 6647
rect 9689 6613 9723 6647
rect 10885 6613 10919 6647
rect 11345 6613 11379 6647
rect 11897 6613 11931 6647
rect 15301 6613 15335 6647
rect 15393 6613 15427 6647
rect 15761 6613 15795 6647
rect 19441 6613 19475 6647
rect 19901 6613 19935 6647
rect 20453 6613 20487 6647
rect 20913 6613 20947 6647
rect 9229 6409 9263 6443
rect 9597 6409 9631 6443
rect 10425 6409 10459 6443
rect 10793 6409 10827 6443
rect 14289 6409 14323 6443
rect 14749 6409 14783 6443
rect 20821 6409 20855 6443
rect 21281 6409 21315 6443
rect 9689 6273 9723 6307
rect 10885 6273 10919 6307
rect 11897 6273 11931 6307
rect 14381 6273 14415 6307
rect 15025 6273 15059 6307
rect 20453 6273 20487 6307
rect 21005 6273 21039 6307
rect 9781 6205 9815 6239
rect 11069 6205 11103 6239
rect 11621 6205 11655 6239
rect 11805 6205 11839 6239
rect 14105 6205 14139 6239
rect 8769 6069 8803 6103
rect 12265 6069 12299 6103
rect 12541 6069 12575 6103
rect 10241 5865 10275 5899
rect 13093 5865 13127 5899
rect 11713 5729 11747 5763
rect 12541 5729 12575 5763
rect 14381 5729 14415 5763
rect 12725 5661 12759 5695
rect 14105 5661 14139 5695
rect 12633 5525 12667 5559
rect 21281 5525 21315 5559
rect 8309 5321 8343 5355
rect 8953 5321 8987 5355
rect 13093 5321 13127 5355
rect 15301 5321 15335 5355
rect 13461 5253 13495 5287
rect 14105 5253 14139 5287
rect 9045 5185 9079 5219
rect 9689 5185 9723 5219
rect 12725 5185 12759 5219
rect 15669 5185 15703 5219
rect 8861 5117 8895 5151
rect 13553 5117 13587 5151
rect 13645 5117 13679 5151
rect 15761 5117 15795 5151
rect 15945 5117 15979 5151
rect 9413 4981 9447 5015
rect 11529 4981 11563 5015
rect 12265 4981 12299 5015
rect 9689 4777 9723 4811
rect 13185 4777 13219 4811
rect 9045 4641 9079 4675
rect 9229 4641 9263 4675
rect 10609 4641 10643 4675
rect 11529 4641 11563 4675
rect 12633 4641 12667 4675
rect 12725 4641 12759 4675
rect 9965 4573 9999 4607
rect 10701 4505 10735 4539
rect 12817 4505 12851 4539
rect 9321 4437 9355 4471
rect 10793 4437 10827 4471
rect 11161 4437 11195 4471
rect 11713 4437 11747 4471
rect 11805 4437 11839 4471
rect 12173 4437 12207 4471
rect 9229 4233 9263 4267
rect 9597 4233 9631 4267
rect 11529 4233 11563 4267
rect 12081 4233 12115 4267
rect 13461 4233 13495 4267
rect 14565 4233 14599 4267
rect 10793 4097 10827 4131
rect 9689 4029 9723 4063
rect 9781 4029 9815 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 13277 4029 13311 4063
rect 13369 4029 13403 4063
rect 14197 4029 14231 4063
rect 11161 3961 11195 3995
rect 13829 3961 13863 3995
rect 15301 3961 15335 3995
rect 14933 3893 14967 3927
rect 15669 3893 15703 3927
rect 9873 3689 9907 3723
rect 10241 3689 10275 3723
rect 10609 3689 10643 3723
rect 11253 3689 11287 3723
rect 15025 3689 15059 3723
rect 16037 3689 16071 3723
rect 17141 3689 17175 3723
rect 14381 3553 14415 3587
rect 14565 3553 14599 3587
rect 15485 3553 15519 3587
rect 16497 3553 16531 3587
rect 16773 3485 16807 3519
rect 14657 3349 14691 3383
rect 15577 3349 15611 3383
rect 15669 3349 15703 3383
rect 15209 3145 15243 3179
rect 15577 3009 15611 3043
rect 16221 2805 16255 2839
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 9677 20587 9735 20593
rect 9677 20553 9689 20587
rect 9723 20584 9735 20587
rect 13078 20584 13084 20596
rect 9723 20556 13084 20584
rect 9723 20553 9735 20556
rect 9677 20547 9735 20553
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 20349 20587 20407 20593
rect 20349 20553 20361 20587
rect 20395 20584 20407 20587
rect 20622 20584 20628 20596
rect 20395 20556 20628 20584
rect 20395 20553 20407 20556
rect 20349 20547 20407 20553
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 20809 20587 20867 20593
rect 20809 20553 20821 20587
rect 20855 20584 20867 20587
rect 21542 20584 21548 20596
rect 20855 20556 21548 20584
rect 20855 20553 20867 20556
rect 20809 20547 20867 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 7282 20476 7288 20528
rect 7340 20516 7346 20528
rect 7340 20488 16574 20516
rect 7340 20476 7346 20488
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10594 20448 10600 20460
rect 9907 20420 10600 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 16546 20448 16574 20488
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16546 20420 16957 20448
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 16945 20411 17003 20417
rect 19904 20420 20637 20448
rect 9306 20340 9312 20392
rect 9364 20380 9370 20392
rect 17310 20380 17316 20392
rect 9364 20352 17316 20380
rect 9364 20340 9370 20352
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 5718 20272 5724 20324
rect 5776 20312 5782 20324
rect 19610 20312 19616 20324
rect 5776 20284 19616 20312
rect 5776 20272 5782 20284
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 17129 20247 17187 20253
rect 17129 20213 17141 20247
rect 17175 20244 17187 20247
rect 18138 20244 18144 20256
rect 17175 20216 18144 20244
rect 17175 20213 17187 20216
rect 17129 20207 17187 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18782 20244 18788 20256
rect 18743 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 19904 20253 19932 20420
rect 20625 20417 20637 20420
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 19889 20247 19947 20253
rect 19889 20244 19901 20247
rect 18932 20216 19901 20244
rect 18932 20204 18938 20216
rect 19889 20213 19901 20216
rect 19935 20213 19947 20247
rect 21174 20244 21180 20256
rect 21135 20216 21180 20244
rect 19889 20207 19947 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 5718 20040 5724 20052
rect 5679 20012 5724 20040
rect 5718 20000 5724 20012
rect 5776 20000 5782 20052
rect 11701 20043 11759 20049
rect 11701 20009 11713 20043
rect 11747 20040 11759 20043
rect 11974 20040 11980 20052
rect 11747 20012 11980 20040
rect 11747 20009 11759 20012
rect 11701 20003 11759 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 17862 20040 17868 20052
rect 12084 20012 17868 20040
rect 7377 19975 7435 19981
rect 7377 19941 7389 19975
rect 7423 19972 7435 19975
rect 12084 19972 12112 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18049 20043 18107 20049
rect 18049 20009 18061 20043
rect 18095 20040 18107 20043
rect 18598 20040 18604 20052
rect 18095 20012 18604 20040
rect 18095 20009 18107 20012
rect 18049 20003 18107 20009
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 19337 20043 19395 20049
rect 19337 20009 19349 20043
rect 19383 20040 19395 20043
rect 20254 20040 20260 20052
rect 19383 20012 20260 20040
rect 19383 20009 19395 20012
rect 19337 20003 19395 20009
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 7423 19944 12112 19972
rect 14829 19975 14887 19981
rect 7423 19941 7435 19944
rect 7377 19935 7435 19941
rect 14829 19941 14841 19975
rect 14875 19972 14887 19975
rect 17497 19975 17555 19981
rect 14875 19944 16574 19972
rect 14875 19941 14887 19944
rect 14829 19935 14887 19941
rect 9122 19904 9128 19916
rect 6886 19876 9128 19904
rect 4154 19836 4160 19848
rect 4115 19808 4160 19836
rect 4154 19796 4160 19808
rect 4212 19796 4218 19848
rect 4706 19836 4712 19848
rect 4667 19808 4712 19836
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19836 5963 19839
rect 6886 19836 6914 19876
rect 9122 19864 9128 19876
rect 9180 19864 9186 19916
rect 9217 19907 9275 19913
rect 9217 19873 9229 19907
rect 9263 19904 9275 19907
rect 9306 19904 9312 19916
rect 9263 19876 9312 19904
rect 9263 19873 9275 19876
rect 9217 19867 9275 19873
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 10413 19907 10471 19913
rect 10413 19873 10425 19907
rect 10459 19904 10471 19907
rect 12250 19904 12256 19916
rect 10459 19876 12256 19904
rect 10459 19873 10471 19876
rect 10413 19867 10471 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 16546 19904 16574 19944
rect 17497 19941 17509 19975
rect 17543 19972 17555 19975
rect 17954 19972 17960 19984
rect 17543 19944 17960 19972
rect 17543 19941 17555 19944
rect 17497 19935 17555 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 18509 19975 18567 19981
rect 18509 19941 18521 19975
rect 18555 19972 18567 19975
rect 19702 19972 19708 19984
rect 18555 19944 19708 19972
rect 18555 19941 18567 19944
rect 18509 19935 18567 19941
rect 19702 19932 19708 19944
rect 19760 19932 19766 19984
rect 19889 19975 19947 19981
rect 19889 19941 19901 19975
rect 19935 19972 19947 19975
rect 20806 19972 20812 19984
rect 19935 19944 20812 19972
rect 19935 19941 19947 19944
rect 19889 19935 19947 19941
rect 20806 19932 20812 19944
rect 20864 19932 20870 19984
rect 19242 19904 19248 19916
rect 16546 19876 19248 19904
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 20993 19907 21051 19913
rect 20993 19873 21005 19907
rect 21039 19904 21051 19907
rect 21266 19904 21272 19916
rect 21039 19876 21272 19904
rect 21039 19873 21051 19876
rect 20993 19867 21051 19873
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 5951 19808 6914 19836
rect 7193 19839 7251 19845
rect 5951 19805 5963 19808
rect 5905 19799 5963 19805
rect 7193 19805 7205 19839
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 9447 19808 9812 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 4985 19771 5043 19777
rect 4985 19737 4997 19771
rect 5031 19768 5043 19771
rect 7208 19768 7236 19799
rect 5031 19740 7236 19768
rect 5031 19737 5043 19740
rect 4985 19731 5043 19737
rect 4338 19700 4344 19712
rect 4299 19672 4344 19700
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 9784 19709 9812 19808
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11517 19839 11575 19845
rect 11517 19836 11529 19839
rect 11296 19808 11529 19836
rect 11296 19796 11302 19808
rect 11517 19805 11529 19808
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 11756 19808 14657 19836
rect 11756 19796 11762 19808
rect 14645 19805 14657 19808
rect 14691 19805 14703 19839
rect 15194 19836 15200 19848
rect 15155 19808 15200 19836
rect 14645 19799 14703 19805
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 16761 19839 16819 19845
rect 16761 19805 16773 19839
rect 16807 19836 16819 19839
rect 17126 19836 17132 19848
rect 16807 19808 17132 19836
rect 16807 19805 16819 19808
rect 16761 19799 16819 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17310 19836 17316 19848
rect 17271 19808 17316 19836
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 17865 19839 17923 19845
rect 17865 19836 17877 19839
rect 17828 19808 17877 19836
rect 17828 19796 17834 19808
rect 17865 19805 17877 19808
rect 17911 19805 17923 19839
rect 17865 19799 17923 19805
rect 18230 19796 18236 19848
rect 18288 19836 18294 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18288 19808 18705 19836
rect 18288 19796 18294 19808
rect 18693 19805 18705 19808
rect 18739 19836 18751 19839
rect 18782 19836 18788 19848
rect 18739 19808 18788 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 19518 19836 19524 19848
rect 19479 19808 19524 19836
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19836 20131 19839
rect 20254 19836 20260 19848
rect 20119 19808 20260 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20254 19796 20260 19808
rect 20312 19796 20318 19848
rect 20622 19796 20628 19848
rect 20680 19836 20686 19848
rect 21177 19839 21235 19845
rect 21177 19836 21189 19839
rect 20680 19808 21189 19836
rect 20680 19796 20686 19808
rect 21177 19805 21189 19808
rect 21223 19805 21235 19839
rect 21177 19799 21235 19805
rect 10137 19771 10195 19777
rect 10137 19737 10149 19771
rect 10183 19768 10195 19771
rect 10781 19771 10839 19777
rect 10781 19768 10793 19771
rect 10183 19740 10793 19768
rect 10183 19737 10195 19740
rect 10137 19731 10195 19737
rect 10781 19737 10793 19740
rect 10827 19737 10839 19771
rect 18414 19768 18420 19780
rect 10781 19731 10839 19737
rect 16546 19740 18420 19768
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19669 9827 19703
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 9769 19663 9827 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 15381 19703 15439 19709
rect 15381 19669 15393 19703
rect 15427 19700 15439 19703
rect 16546 19700 16574 19740
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 15427 19672 16574 19700
rect 16945 19703 17003 19709
rect 15427 19669 15439 19672
rect 15381 19663 15439 19669
rect 16945 19669 16957 19703
rect 16991 19700 17003 19703
rect 17678 19700 17684 19712
rect 16991 19672 17684 19700
rect 16991 19669 17003 19672
rect 16945 19663 17003 19669
rect 17678 19660 17684 19672
rect 17736 19660 17742 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 3878 19496 3884 19508
rect 3839 19468 3884 19496
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 9861 19499 9919 19505
rect 9861 19465 9873 19499
rect 9907 19496 9919 19499
rect 13722 19496 13728 19508
rect 9907 19468 13728 19496
rect 9907 19465 9919 19468
rect 9861 19459 9919 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 21358 19496 21364 19508
rect 20763 19468 21364 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 1394 19388 1400 19440
rect 1452 19428 1458 19440
rect 2590 19428 2596 19440
rect 1452 19400 2596 19428
rect 1452 19388 1458 19400
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 4246 19388 4252 19440
rect 4304 19428 4310 19440
rect 4798 19428 4804 19440
rect 4304 19400 4804 19428
rect 4304 19388 4310 19400
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 7282 19428 7288 19440
rect 7243 19400 7288 19428
rect 7282 19388 7288 19400
rect 7340 19388 7346 19440
rect 10689 19431 10747 19437
rect 10060 19400 10640 19428
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4522 19360 4528 19372
rect 4111 19332 4528 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 4522 19320 4528 19332
rect 4580 19320 4586 19372
rect 7558 19360 7564 19372
rect 7519 19332 7564 19360
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 10060 19369 10088 19400
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19329 10103 19363
rect 10410 19360 10416 19372
rect 10371 19332 10416 19360
rect 10045 19323 10103 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 10612 19360 10640 19400
rect 10689 19397 10701 19431
rect 10735 19428 10747 19431
rect 11698 19428 11704 19440
rect 10735 19400 11704 19428
rect 10735 19397 10747 19400
rect 10689 19391 10747 19397
rect 11698 19388 11704 19400
rect 11756 19388 11762 19440
rect 12652 19431 12710 19437
rect 12652 19397 12664 19431
rect 12698 19428 12710 19431
rect 12894 19428 12900 19440
rect 12698 19400 12900 19428
rect 12698 19397 12710 19400
rect 12652 19391 12710 19397
rect 12894 19388 12900 19400
rect 12952 19388 12958 19440
rect 15378 19388 15384 19440
rect 15436 19428 15442 19440
rect 16390 19428 16396 19440
rect 15436 19400 16396 19428
rect 15436 19388 15442 19400
rect 16390 19388 16396 19400
rect 16448 19388 16454 19440
rect 17862 19428 17868 19440
rect 17328 19400 17868 19428
rect 10778 19360 10784 19372
rect 10612 19332 10784 19360
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 14366 19360 14372 19372
rect 11572 19332 14372 19360
rect 11572 19320 11578 19332
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 17328 19369 17356 19400
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 20990 19388 20996 19440
rect 21048 19428 21054 19440
rect 22462 19428 22468 19440
rect 21048 19400 22468 19428
rect 21048 19388 21054 19400
rect 22462 19388 22468 19400
rect 22520 19388 22526 19440
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17569 19363 17627 19369
rect 17569 19360 17581 19363
rect 17313 19323 17371 19329
rect 17420 19332 17581 19360
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 6638 19292 6644 19304
rect 4028 19264 6644 19292
rect 4028 19252 4034 19264
rect 6638 19252 6644 19264
rect 6696 19252 6702 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 10870 19292 10876 19304
rect 9824 19264 10876 19292
rect 9824 19252 9830 19264
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 13262 19292 13268 19304
rect 12943 19264 13268 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 16942 19252 16948 19304
rect 17000 19292 17006 19304
rect 17420 19292 17448 19332
rect 17569 19329 17581 19332
rect 17615 19329 17627 19363
rect 17569 19323 17627 19329
rect 18506 19320 18512 19372
rect 18564 19360 18570 19372
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 18564 19332 20913 19360
rect 18564 19320 18570 19332
rect 20901 19329 20913 19332
rect 20947 19360 20959 19363
rect 21174 19360 21180 19372
rect 20947 19332 21180 19360
rect 20947 19329 20959 19332
rect 20901 19323 20959 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 17000 19264 17448 19292
rect 17000 19252 17006 19264
rect 934 19184 940 19236
rect 992 19224 998 19236
rect 5810 19224 5816 19236
rect 992 19196 5816 19224
rect 992 19184 998 19196
rect 5810 19184 5816 19196
rect 5868 19184 5874 19236
rect 6886 19196 11652 19224
rect 4338 19116 4344 19168
rect 4396 19156 4402 19168
rect 6886 19156 6914 19196
rect 11514 19156 11520 19168
rect 4396 19128 6914 19156
rect 11475 19128 11520 19156
rect 4396 19116 4402 19128
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11624 19156 11652 19196
rect 12912 19196 16574 19224
rect 12912 19156 12940 19196
rect 13262 19156 13268 19168
rect 11624 19128 12940 19156
rect 13175 19128 13268 19156
rect 13262 19116 13268 19128
rect 13320 19156 13326 19168
rect 13722 19156 13728 19168
rect 13320 19128 13728 19156
rect 13320 19116 13326 19128
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 16546 19156 16574 19196
rect 19518 19184 19524 19236
rect 19576 19224 19582 19236
rect 19705 19227 19763 19233
rect 19705 19224 19717 19227
rect 19576 19196 19717 19224
rect 19576 19184 19582 19196
rect 19705 19193 19717 19196
rect 19751 19224 19763 19227
rect 20438 19224 20444 19236
rect 19751 19196 20444 19224
rect 19751 19193 19763 19196
rect 19705 19187 19763 19193
rect 20438 19184 20444 19196
rect 20496 19184 20502 19236
rect 18598 19156 18604 19168
rect 16546 19128 18604 19156
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 18690 19116 18696 19168
rect 18748 19156 18754 19168
rect 19058 19156 19064 19168
rect 18748 19128 18793 19156
rect 19019 19128 19064 19156
rect 18748 19116 18754 19128
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 20254 19156 20260 19168
rect 20215 19128 20260 19156
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 7374 18952 7380 18964
rect 3200 18924 7380 18952
rect 3200 18912 3206 18924
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 16298 18952 16304 18964
rect 8496 18924 16304 18952
rect 4080 18856 8248 18884
rect 4080 18825 4108 18856
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 2406 18748 2412 18760
rect 2367 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 5166 18748 5172 18760
rect 4295 18720 5028 18748
rect 5127 18720 5172 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 2133 18683 2191 18689
rect 2133 18649 2145 18683
rect 2179 18680 2191 18683
rect 4154 18680 4160 18692
rect 2179 18652 4160 18680
rect 2179 18649 2191 18652
rect 2133 18643 2191 18649
rect 4154 18640 4160 18652
rect 4212 18640 4218 18692
rect 4890 18680 4896 18692
rect 4851 18652 4896 18680
rect 4890 18640 4896 18652
rect 4948 18640 4954 18692
rect 5000 18680 5028 18720
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 7742 18680 7748 18692
rect 5000 18652 7748 18680
rect 7742 18640 7748 18652
rect 7800 18640 7806 18692
rect 8220 18680 8248 18856
rect 8496 18825 8524 18924
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18785 8539 18819
rect 9122 18816 9128 18828
rect 9083 18788 9128 18816
rect 8481 18779 8539 18785
rect 9122 18776 9128 18788
rect 9180 18776 9186 18828
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 8662 18748 8668 18760
rect 8343 18720 8668 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 8941 18751 8999 18757
rect 8941 18717 8953 18751
rect 8987 18748 8999 18751
rect 9030 18748 9036 18760
rect 8987 18720 9036 18748
rect 8987 18717 8999 18720
rect 8941 18711 8999 18717
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 12115 18720 12357 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12345 18717 12357 18720
rect 12391 18748 12403 18751
rect 12434 18748 12440 18760
rect 12391 18720 12440 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 12434 18708 12440 18720
rect 12492 18748 12498 18760
rect 13722 18748 13728 18760
rect 12492 18720 13728 18748
rect 12492 18708 12498 18720
rect 13722 18708 13728 18720
rect 13780 18748 13786 18760
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 13780 18720 14197 18748
rect 13780 18708 13786 18720
rect 14185 18717 14197 18720
rect 14231 18748 14243 18751
rect 14921 18751 14979 18757
rect 14921 18748 14933 18751
rect 14231 18720 14933 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14921 18717 14933 18720
rect 14967 18748 14979 18751
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 14967 18720 16681 18748
rect 14967 18717 14979 18720
rect 14921 18711 14979 18717
rect 16669 18717 16681 18720
rect 16715 18748 16727 18751
rect 17862 18748 17868 18760
rect 16715 18720 17868 18748
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 17862 18708 17868 18720
rect 17920 18748 17926 18760
rect 18693 18751 18751 18757
rect 18693 18748 18705 18751
rect 17920 18720 18705 18748
rect 17920 18708 17926 18720
rect 18693 18717 18705 18720
rect 18739 18748 18751 18751
rect 19058 18748 19064 18760
rect 18739 18720 19064 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 19058 18708 19064 18720
rect 19116 18748 19122 18760
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 19116 18720 19349 18748
rect 19116 18708 19122 18720
rect 19337 18717 19349 18720
rect 19383 18748 19395 18751
rect 19889 18751 19947 18757
rect 19889 18748 19901 18751
rect 19383 18720 19901 18748
rect 19383 18717 19395 18720
rect 19337 18711 19395 18717
rect 19889 18717 19901 18720
rect 19935 18748 19947 18751
rect 21266 18748 21272 18760
rect 19935 18720 21272 18748
rect 19935 18717 19947 18720
rect 19889 18711 19947 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 11054 18680 11060 18692
rect 8220 18652 11060 18680
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 11146 18640 11152 18692
rect 11204 18680 11210 18692
rect 11802 18683 11860 18689
rect 11802 18680 11814 18683
rect 11204 18652 11814 18680
rect 11204 18640 11210 18652
rect 11802 18649 11814 18652
rect 11848 18680 11860 18683
rect 11974 18680 11980 18692
rect 11848 18652 11980 18680
rect 11848 18649 11860 18652
rect 11802 18643 11860 18649
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 12612 18683 12670 18689
rect 12612 18649 12624 18683
rect 12658 18680 12670 18683
rect 13170 18680 13176 18692
rect 12658 18652 13176 18680
rect 12658 18649 12670 18652
rect 12612 18643 12670 18649
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 15188 18683 15246 18689
rect 13280 18652 13860 18680
rect 7834 18612 7840 18624
rect 7795 18584 7840 18612
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 8202 18612 8208 18624
rect 8115 18584 8208 18612
rect 8202 18572 8208 18584
rect 8260 18612 8266 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 8260 18584 9689 18612
rect 8260 18572 8266 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 10686 18612 10692 18624
rect 10647 18584 10692 18612
rect 9677 18575 9735 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 13280 18612 13308 18652
rect 11756 18584 13308 18612
rect 11756 18572 11762 18584
rect 13630 18572 13636 18624
rect 13688 18612 13694 18624
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13688 18584 13737 18612
rect 13688 18572 13694 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 13832 18612 13860 18652
rect 15188 18649 15200 18683
rect 15234 18680 15246 18683
rect 15470 18680 15476 18692
rect 15234 18652 15476 18680
rect 15234 18649 15246 18652
rect 15188 18643 15246 18649
rect 15470 18640 15476 18652
rect 15528 18640 15534 18692
rect 17126 18680 17132 18692
rect 15580 18652 17132 18680
rect 15580 18612 15608 18652
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 17494 18640 17500 18692
rect 17552 18680 17558 18692
rect 18426 18683 18484 18689
rect 18426 18680 18438 18683
rect 17552 18652 18438 18680
rect 17552 18640 17558 18652
rect 18426 18649 18438 18652
rect 18472 18649 18484 18683
rect 18426 18643 18484 18649
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 20134 18683 20192 18689
rect 20134 18680 20146 18683
rect 19576 18652 20146 18680
rect 19576 18640 19582 18652
rect 20134 18649 20146 18652
rect 20180 18649 20192 18683
rect 20134 18643 20192 18649
rect 13832 18584 15608 18612
rect 13725 18575 13783 18581
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 16942 18612 16948 18624
rect 16356 18584 16948 18612
rect 16356 18572 16362 18584
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17310 18612 17316 18624
rect 17271 18584 17316 18612
rect 17310 18572 17316 18584
rect 17368 18572 17374 18624
rect 21174 18572 21180 18624
rect 21232 18612 21238 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 21232 18584 21281 18612
rect 21232 18572 21238 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 382 18368 388 18420
rect 440 18408 446 18420
rect 6454 18408 6460 18420
rect 440 18380 6460 18408
rect 440 18368 446 18380
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 8662 18408 8668 18420
rect 8623 18380 8668 18408
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 12069 18411 12127 18417
rect 12069 18377 12081 18411
rect 12115 18408 12127 18411
rect 12434 18408 12440 18420
rect 12115 18380 12440 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 12710 18408 12716 18420
rect 12584 18380 12716 18408
rect 12584 18368 12590 18380
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 14001 18411 14059 18417
rect 14001 18408 14013 18411
rect 13780 18380 14013 18408
rect 13780 18368 13786 18380
rect 14001 18377 14013 18380
rect 14047 18377 14059 18411
rect 14001 18371 14059 18377
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 17402 18408 17408 18420
rect 17000 18380 17408 18408
rect 17000 18368 17006 18380
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 20625 18411 20683 18417
rect 20625 18408 20637 18411
rect 19024 18380 20637 18408
rect 19024 18368 19030 18380
rect 20625 18377 20637 18380
rect 20671 18377 20683 18411
rect 20625 18371 20683 18377
rect 4522 18340 4528 18352
rect 4483 18312 4528 18340
rect 4522 18300 4528 18312
rect 4580 18300 4586 18352
rect 10686 18340 10692 18352
rect 6656 18312 10692 18340
rect 4798 18272 4804 18284
rect 4759 18244 4804 18272
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 6656 18213 6684 18312
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 11054 18300 11060 18352
rect 11112 18340 11118 18352
rect 15194 18340 15200 18352
rect 11112 18312 15200 18340
rect 11112 18300 11118 18312
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 20898 18340 20904 18352
rect 16546 18312 20904 18340
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 7561 18275 7619 18281
rect 7561 18272 7573 18275
rect 6963 18244 7573 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 7561 18241 7573 18244
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 8662 18272 8668 18284
rect 7800 18244 8668 18272
rect 7800 18232 7806 18244
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18272 9459 18275
rect 10045 18275 10103 18281
rect 10045 18272 10057 18275
rect 9447 18244 10057 18272
rect 9447 18241 9459 18244
rect 9401 18235 9459 18241
rect 10045 18241 10057 18244
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 13458 18275 13516 18281
rect 13458 18272 13470 18275
rect 11020 18244 13470 18272
rect 11020 18232 11026 18244
rect 13458 18241 13470 18244
rect 13504 18272 13516 18275
rect 13630 18272 13636 18284
rect 13504 18244 13636 18272
rect 13504 18241 13516 18244
rect 13458 18235 13516 18241
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 13780 18244 13825 18272
rect 13780 18232 13786 18244
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18173 6699 18207
rect 6822 18204 6828 18216
rect 6783 18176 6828 18204
rect 6641 18167 6699 18173
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 9364 18176 9505 18204
rect 9364 18164 9370 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18204 9643 18207
rect 16546 18204 16574 18312
rect 20898 18300 20904 18312
rect 20956 18340 20962 18352
rect 21174 18340 21180 18352
rect 20956 18312 21180 18340
rect 20956 18300 20962 18312
rect 21174 18300 21180 18312
rect 21232 18300 21238 18352
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18305 18275 18363 18281
rect 18305 18272 18317 18275
rect 18196 18244 18317 18272
rect 18196 18232 18202 18244
rect 18305 18241 18317 18244
rect 18351 18272 18363 18275
rect 18690 18272 18696 18284
rect 18351 18244 18696 18272
rect 18351 18241 18363 18244
rect 18305 18235 18363 18241
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18272 20315 18275
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20303 18244 20821 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 20809 18241 20821 18244
rect 20855 18272 20867 18275
rect 21450 18272 21456 18284
rect 20855 18244 21456 18272
rect 20855 18241 20867 18244
rect 20809 18235 20867 18241
rect 21450 18232 21456 18244
rect 21508 18232 21514 18284
rect 9631 18176 12756 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 4890 18096 4896 18148
rect 4948 18136 4954 18148
rect 11698 18136 11704 18148
rect 4948 18108 11704 18136
rect 4948 18096 4954 18108
rect 11698 18096 11704 18108
rect 11756 18096 11762 18148
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 6914 18068 6920 18080
rect 6604 18040 6920 18068
rect 6604 18028 6610 18040
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 7282 18068 7288 18080
rect 7243 18040 7288 18068
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 9490 18028 9496 18080
rect 9548 18068 9554 18080
rect 12342 18068 12348 18080
rect 9548 18040 12348 18068
rect 9548 18028 9554 18040
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 12728 18068 12756 18176
rect 13740 18176 16574 18204
rect 13740 18068 13768 18176
rect 17862 18164 17868 18216
rect 17920 18204 17926 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17920 18176 18061 18204
rect 17920 18164 17926 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 14274 18096 14280 18148
rect 14332 18136 14338 18148
rect 17494 18136 17500 18148
rect 14332 18108 17500 18136
rect 14332 18096 14338 18108
rect 17494 18096 17500 18108
rect 17552 18096 17558 18148
rect 19797 18139 19855 18145
rect 19797 18105 19809 18139
rect 19843 18136 19855 18139
rect 19843 18108 21312 18136
rect 19843 18105 19855 18108
rect 19797 18099 19855 18105
rect 21284 18080 21312 18108
rect 12728 18040 13768 18068
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 15286 18068 15292 18080
rect 13872 18040 15292 18068
rect 13872 18028 13878 18040
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 19518 18068 19524 18080
rect 19475 18040 19524 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 21266 18068 21272 18080
rect 21227 18040 21272 18068
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 4706 17864 4712 17876
rect 4571 17836 4712 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 9769 17867 9827 17873
rect 5960 17836 9720 17864
rect 5960 17824 5966 17836
rect 6457 17799 6515 17805
rect 6457 17796 6469 17799
rect 5460 17768 6469 17796
rect 3878 17728 3884 17740
rect 3839 17700 3884 17728
rect 3878 17688 3884 17700
rect 3936 17688 3942 17740
rect 5460 17737 5488 17768
rect 6457 17765 6469 17768
rect 6503 17796 6515 17799
rect 9582 17796 9588 17808
rect 6503 17768 9588 17796
rect 6503 17765 6515 17768
rect 6457 17759 6515 17765
rect 9582 17756 9588 17768
rect 9640 17756 9646 17808
rect 9692 17796 9720 17836
rect 9769 17833 9781 17867
rect 9815 17864 9827 17867
rect 10226 17864 10232 17876
rect 9815 17836 10232 17864
rect 9815 17833 9827 17836
rect 9769 17827 9827 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 13170 17864 13176 17876
rect 10336 17836 12848 17864
rect 13131 17836 13176 17864
rect 10336 17796 10364 17836
rect 9692 17768 10364 17796
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17697 5503 17731
rect 5626 17728 5632 17740
rect 5587 17700 5632 17728
rect 5445 17691 5503 17697
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 9214 17728 9220 17740
rect 5736 17700 9076 17728
rect 9175 17700 9220 17728
rect 3896 17660 3924 17688
rect 5736 17660 5764 17700
rect 3896 17632 5764 17660
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 9048 17660 9076 17700
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 9309 17731 9367 17737
rect 9309 17697 9321 17731
rect 9355 17728 9367 17731
rect 10318 17728 10324 17740
rect 9355 17700 10324 17728
rect 9355 17697 9367 17700
rect 9309 17691 9367 17697
rect 10318 17688 10324 17700
rect 10376 17728 10382 17740
rect 10413 17731 10471 17737
rect 10413 17728 10425 17731
rect 10376 17700 10425 17728
rect 10376 17688 10382 17700
rect 10413 17697 10425 17700
rect 10459 17697 10471 17731
rect 10413 17691 10471 17697
rect 11793 17663 11851 17669
rect 6052 17632 8432 17660
rect 9048 17632 10640 17660
rect 6052 17620 6058 17632
rect 4065 17595 4123 17601
rect 4065 17561 4077 17595
rect 4111 17592 4123 17595
rect 5353 17595 5411 17601
rect 4111 17564 5028 17592
rect 4111 17561 4123 17564
rect 4065 17555 4123 17561
rect 4157 17527 4215 17533
rect 4157 17493 4169 17527
rect 4203 17524 4215 17527
rect 4338 17524 4344 17536
rect 4203 17496 4344 17524
rect 4203 17493 4215 17496
rect 4157 17487 4215 17493
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 5000 17533 5028 17564
rect 5353 17561 5365 17595
rect 5399 17592 5411 17595
rect 6089 17595 6147 17601
rect 6089 17592 6101 17595
rect 5399 17564 6101 17592
rect 5399 17561 5411 17564
rect 5353 17555 5411 17561
rect 6089 17561 6101 17564
rect 6135 17592 6147 17595
rect 7190 17592 7196 17604
rect 6135 17564 7196 17592
rect 6135 17561 6147 17564
rect 6089 17555 6147 17561
rect 7190 17552 7196 17564
rect 7248 17552 7254 17604
rect 4985 17527 5043 17533
rect 4985 17493 4997 17527
rect 5031 17493 5043 17527
rect 8404 17524 8432 17632
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 8536 17564 9413 17592
rect 8536 17552 8542 17564
rect 9401 17561 9413 17564
rect 9447 17592 9459 17595
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 9447 17564 10057 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 10045 17561 10057 17564
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 9582 17524 9588 17536
rect 8404 17496 9588 17524
rect 4985 17487 5043 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10502 17524 10508 17536
rect 9732 17496 10508 17524
rect 9732 17484 9738 17496
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 10612 17524 10640 17632
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 12434 17660 12440 17672
rect 11839 17632 12440 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 10686 17552 10692 17604
rect 10744 17592 10750 17604
rect 12038 17595 12096 17601
rect 12038 17592 12050 17595
rect 10744 17564 12050 17592
rect 10744 17552 10750 17564
rect 12038 17561 12050 17564
rect 12084 17561 12096 17595
rect 12820 17592 12848 17836
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 13541 17867 13599 17873
rect 13541 17833 13553 17867
rect 13587 17864 13599 17867
rect 13722 17864 13728 17876
rect 13587 17836 13728 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 17221 17867 17279 17873
rect 17221 17833 17233 17867
rect 17267 17864 17279 17867
rect 17862 17864 17868 17876
rect 17267 17836 17868 17864
rect 17267 17833 17279 17836
rect 17221 17827 17279 17833
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17236 17728 17264 17827
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 16899 17700 17264 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 16597 17663 16655 17669
rect 16597 17660 16609 17663
rect 13136 17632 16609 17660
rect 13136 17620 13142 17632
rect 16597 17629 16609 17632
rect 16643 17660 16655 17663
rect 17310 17660 17316 17672
rect 16643 17632 17316 17660
rect 16643 17629 16655 17632
rect 16597 17623 16655 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 20898 17620 20904 17672
rect 20956 17669 20962 17672
rect 20956 17660 20968 17669
rect 21177 17663 21235 17669
rect 20956 17632 21001 17660
rect 20956 17623 20968 17632
rect 21177 17629 21189 17663
rect 21223 17660 21235 17663
rect 21266 17660 21272 17672
rect 21223 17632 21272 17660
rect 21223 17629 21235 17632
rect 21177 17623 21235 17629
rect 20956 17620 20962 17623
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 18138 17592 18144 17604
rect 12820 17564 18144 17592
rect 12038 17555 12096 17561
rect 18138 17552 18144 17564
rect 18196 17552 18202 17604
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 10612 17496 15485 17524
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 19797 17527 19855 17533
rect 19797 17524 19809 17527
rect 19760 17496 19809 17524
rect 19760 17484 19766 17496
rect 19797 17493 19809 17496
rect 19843 17493 19855 17527
rect 19797 17487 19855 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 4338 17320 4344 17332
rect 4299 17292 4344 17320
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 4856 17292 5273 17320
rect 4856 17280 4862 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 5626 17280 5632 17332
rect 5684 17320 5690 17332
rect 10229 17323 10287 17329
rect 5684 17292 9536 17320
rect 5684 17280 5690 17292
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 7834 17252 7840 17264
rect 5767 17224 7840 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 5675 17156 6377 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 6972 17156 7017 17184
rect 6972 17144 6978 17156
rect 5902 17116 5908 17128
rect 5863 17088 5908 17116
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 9508 16980 9536 17292
rect 10229 17289 10241 17323
rect 10275 17320 10287 17323
rect 10410 17320 10416 17332
rect 10275 17292 10416 17320
rect 10275 17289 10287 17292
rect 10229 17283 10287 17289
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 10612 17292 16574 17320
rect 10612 17252 10640 17292
rect 12434 17252 12440 17264
rect 9692 17224 10640 17252
rect 11532 17224 12440 17252
rect 9692 17184 9720 17224
rect 11532 17193 11560 17224
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 15746 17252 15752 17264
rect 14108 17224 15752 17252
rect 9600 17156 9720 17184
rect 9861 17187 9919 17193
rect 9600 17125 9628 17156
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 9907 17156 10517 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 10505 17153 10517 17156
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 11606 17184 11612 17196
rect 11563 17156 11612 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 11790 17193 11796 17196
rect 11784 17147 11796 17193
rect 11848 17184 11854 17196
rect 11848 17156 11884 17184
rect 11790 17144 11796 17147
rect 11848 17144 11854 17156
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12400 17156 13216 17184
rect 12400 17144 12406 17156
rect 9585 17119 9643 17125
rect 9585 17085 9597 17119
rect 9631 17085 9643 17119
rect 9766 17116 9772 17128
rect 9727 17088 9772 17116
rect 9585 17079 9643 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 11146 17048 11152 17060
rect 9732 17020 11152 17048
rect 9732 17008 9738 17020
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 13078 17048 13084 17060
rect 12452 17020 13084 17048
rect 12452 16980 12480 17020
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 9508 16952 12480 16980
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 12986 16980 12992 16992
rect 12943 16952 12992 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13188 16980 13216 17156
rect 14108 17125 14136 17224
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 14366 17193 14372 17196
rect 14360 17184 14372 17193
rect 14327 17156 14372 17184
rect 14360 17147 14372 17156
rect 14366 17144 14372 17147
rect 14424 17144 14430 17196
rect 16546 17184 16574 17292
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 18325 17323 18383 17329
rect 18325 17320 18337 17323
rect 17920 17292 18337 17320
rect 17920 17280 17926 17292
rect 18064 17193 18092 17292
rect 18325 17289 18337 17292
rect 18371 17289 18383 17323
rect 18325 17283 18383 17289
rect 17793 17187 17851 17193
rect 17793 17184 17805 17187
rect 16546 17156 17805 17184
rect 17793 17153 17805 17156
rect 17839 17184 17851 17187
rect 18049 17187 18107 17193
rect 17839 17156 18000 17184
rect 17839 17153 17851 17156
rect 17793 17147 17851 17153
rect 13265 17119 13323 17125
rect 13265 17085 13277 17119
rect 13311 17116 13323 17119
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13311 17088 14105 17116
rect 13311 17085 13323 17088
rect 13265 17079 13323 17085
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 17972 17116 18000 17156
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 19702 17144 19708 17196
rect 19760 17184 19766 17196
rect 20634 17187 20692 17193
rect 20634 17184 20646 17187
rect 19760 17156 20646 17184
rect 19760 17144 19766 17156
rect 20634 17153 20646 17156
rect 20680 17153 20692 17187
rect 20634 17147 20692 17153
rect 20901 17119 20959 17125
rect 17972 17088 19564 17116
rect 14093 17079 14151 17085
rect 19536 17057 19564 17088
rect 20901 17085 20913 17119
rect 20947 17116 20959 17119
rect 20947 17088 21312 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 15212 17020 16681 17048
rect 15212 16992 15240 17020
rect 16669 17017 16681 17020
rect 16715 17017 16727 17051
rect 16669 17011 16727 17017
rect 19521 17051 19579 17057
rect 19521 17017 19533 17051
rect 19567 17017 19579 17051
rect 19521 17011 19579 17017
rect 21284 16992 21312 17088
rect 15194 16980 15200 16992
rect 13188 16952 15200 16980
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 15470 16980 15476 16992
rect 15431 16952 15476 16980
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 6822 16776 6828 16788
rect 6595 16748 6828 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 6972 16748 7328 16776
rect 6972 16736 6978 16748
rect 4724 16680 7236 16708
rect 4522 16640 4528 16652
rect 4483 16612 4528 16640
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 4724 16649 4752 16680
rect 4709 16643 4767 16649
rect 4709 16609 4721 16643
rect 4755 16609 4767 16643
rect 5994 16640 6000 16652
rect 5955 16612 6000 16640
rect 4709 16603 4767 16609
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 7208 16572 7236 16680
rect 7300 16649 7328 16748
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 12342 16776 12348 16788
rect 9272 16748 12348 16776
rect 9272 16736 9278 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 15470 16776 15476 16788
rect 12636 16748 15476 16776
rect 7392 16680 11468 16708
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 7392 16572 7420 16680
rect 7469 16643 7527 16649
rect 7469 16609 7481 16643
rect 7515 16640 7527 16643
rect 9490 16640 9496 16652
rect 7515 16612 9496 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16640 10287 16643
rect 10962 16640 10968 16652
rect 10275 16612 10968 16640
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11440 16572 11468 16680
rect 11606 16640 11612 16652
rect 11567 16612 11612 16640
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12636 16572 12664 16748
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 20898 16776 20904 16788
rect 20859 16748 20904 16776
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16640 17739 16643
rect 17862 16640 17868 16652
rect 17727 16612 17868 16640
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 15194 16572 15200 16584
rect 15252 16581 15258 16584
rect 7208 16544 7420 16572
rect 7484 16544 10732 16572
rect 11440 16544 12664 16572
rect 15164 16544 15200 16572
rect 5994 16464 6000 16516
rect 6052 16504 6058 16516
rect 6181 16507 6239 16513
rect 6181 16504 6193 16507
rect 6052 16476 6193 16504
rect 6052 16464 6058 16476
rect 6181 16473 6193 16476
rect 6227 16473 6239 16507
rect 6181 16467 6239 16473
rect 7282 16464 7288 16516
rect 7340 16504 7346 16516
rect 7484 16504 7512 16544
rect 7340 16476 7512 16504
rect 9953 16507 10011 16513
rect 7340 16464 7346 16476
rect 9953 16473 9965 16507
rect 9999 16504 10011 16507
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 9999 16476 10609 16504
rect 9999 16473 10011 16476
rect 9953 16467 10011 16473
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 10597 16467 10655 16473
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 4065 16439 4123 16445
rect 4065 16436 4077 16439
rect 2464 16408 4077 16436
rect 2464 16396 2470 16408
rect 4065 16405 4077 16408
rect 4111 16405 4123 16439
rect 4065 16399 4123 16405
rect 4433 16439 4491 16445
rect 4433 16405 4445 16439
rect 4479 16436 4491 16439
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 4479 16408 5089 16436
rect 4479 16405 4491 16408
rect 4433 16399 4491 16405
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 6089 16439 6147 16445
rect 6089 16436 6101 16439
rect 5592 16408 6101 16436
rect 5592 16396 5598 16408
rect 6089 16405 6101 16408
rect 6135 16405 6147 16439
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 6089 16399 6147 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 7190 16396 7196 16448
rect 7248 16436 7254 16448
rect 7834 16436 7840 16448
rect 7248 16408 7840 16436
rect 7248 16396 7254 16408
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 9585 16439 9643 16445
rect 9585 16436 9597 16439
rect 8720 16408 9597 16436
rect 8720 16396 8726 16408
rect 9585 16405 9597 16408
rect 9631 16405 9643 16439
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 9585 16399 9643 16405
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10704 16436 10732 16544
rect 15194 16532 15200 16544
rect 15252 16535 15264 16581
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15746 16572 15752 16584
rect 15519 16544 15752 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15252 16532 15258 16535
rect 15746 16532 15752 16544
rect 15804 16572 15810 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15804 16544 15853 16572
rect 15804 16532 15810 16544
rect 15841 16541 15853 16544
rect 15887 16572 15899 16575
rect 17696 16572 17724 16603
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 21266 16640 21272 16652
rect 21227 16612 21272 16640
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 15887 16544 17724 16572
rect 18233 16575 18291 16581
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16572 18567 16575
rect 20717 16575 20775 16581
rect 20717 16572 20729 16575
rect 18555 16544 20729 16572
rect 18555 16541 18567 16544
rect 18509 16535 18567 16541
rect 20717 16541 20729 16544
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 11698 16464 11704 16516
rect 11756 16504 11762 16516
rect 11854 16507 11912 16513
rect 11854 16504 11866 16507
rect 11756 16476 11866 16504
rect 11756 16464 11762 16476
rect 11854 16473 11866 16476
rect 11900 16473 11912 16507
rect 11854 16467 11912 16473
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 17414 16507 17472 16513
rect 17414 16504 17426 16507
rect 15344 16476 17426 16504
rect 15344 16464 15350 16476
rect 17414 16473 17426 16476
rect 17460 16473 17472 16507
rect 17414 16467 17472 16473
rect 17586 16464 17592 16516
rect 17644 16504 17650 16516
rect 18248 16504 18276 16535
rect 17644 16476 18276 16504
rect 17644 16464 17650 16476
rect 12066 16436 12072 16448
rect 10704 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 12894 16436 12900 16448
rect 12584 16408 12900 16436
rect 12584 16396 12590 16408
rect 12894 16396 12900 16408
rect 12952 16436 12958 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12952 16408 13001 16436
rect 12952 16396 12958 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 13446 16436 13452 16448
rect 13403 16408 13452 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14093 16439 14151 16445
rect 14093 16436 14105 16439
rect 13872 16408 14105 16436
rect 13872 16396 13878 16408
rect 14093 16405 14105 16408
rect 14139 16405 14151 16439
rect 14093 16399 14151 16405
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 16301 16439 16359 16445
rect 16301 16436 16313 16439
rect 15252 16408 16313 16436
rect 15252 16396 15258 16408
rect 16301 16405 16313 16408
rect 16347 16405 16359 16439
rect 16301 16399 16359 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 5592 16204 5641 16232
rect 5592 16192 5598 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 5629 16195 5687 16201
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 8205 16235 8263 16241
rect 5776 16204 6914 16232
rect 5776 16192 5782 16204
rect 5994 16124 6000 16176
rect 6052 16164 6058 16176
rect 6641 16167 6699 16173
rect 6641 16164 6653 16167
rect 6052 16136 6653 16164
rect 6052 16124 6058 16136
rect 6641 16133 6653 16136
rect 6687 16164 6699 16167
rect 6730 16164 6736 16176
rect 6687 16136 6736 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 6886 16096 6914 16204
rect 8205 16201 8217 16235
rect 8251 16232 8263 16235
rect 10042 16232 10048 16244
rect 8251 16204 10048 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 11974 16232 11980 16244
rect 11931 16204 11980 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 17586 16232 17592 16244
rect 12124 16204 17592 16232
rect 12124 16192 12130 16204
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 13170 16164 13176 16176
rect 10336 16136 13176 16164
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6886 16068 7205 16096
rect 7193 16065 7205 16068
rect 7239 16096 7251 16099
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7239 16068 7757 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 7837 16099 7895 16105
rect 7837 16065 7849 16099
rect 7883 16096 7895 16099
rect 8386 16096 8392 16108
rect 7883 16068 8392 16096
rect 7883 16065 7895 16068
rect 7837 16059 7895 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 10336 16028 10364 16136
rect 13170 16124 13176 16136
rect 13228 16124 13234 16176
rect 12986 16056 12992 16108
rect 13044 16105 13050 16108
rect 13044 16096 13056 16105
rect 13044 16068 13089 16096
rect 13044 16059 13056 16068
rect 13044 16056 13050 16059
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 21094 16099 21152 16105
rect 21094 16096 21106 16099
rect 20588 16068 21106 16096
rect 20588 16056 20594 16068
rect 21094 16065 21106 16068
rect 21140 16065 21152 16099
rect 21094 16059 21152 16065
rect 21266 16056 21272 16108
rect 21324 16096 21330 16108
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 21324 16068 21373 16096
rect 21324 16056 21330 16068
rect 21361 16065 21373 16068
rect 21407 16065 21419 16099
rect 21361 16059 21419 16065
rect 7699 16000 10364 16028
rect 13265 16031 13323 16037
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 13311 16000 13492 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 13464 15904 13492 16000
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8481 15895 8539 15901
rect 8481 15892 8493 15895
rect 8444 15864 8493 15892
rect 8444 15852 8450 15864
rect 8481 15861 8493 15864
rect 8527 15861 8539 15895
rect 8481 15855 8539 15861
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 13504 15864 13553 15892
rect 13504 15852 13510 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 19058 15892 19064 15904
rect 14516 15864 19064 15892
rect 14516 15852 14522 15864
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 19978 15892 19984 15904
rect 19939 15864 19984 15892
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 19337 15691 19395 15697
rect 19337 15657 19349 15691
rect 19383 15688 19395 15691
rect 21266 15688 21272 15700
rect 19383 15660 21272 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 14274 15552 14280 15564
rect 13188 15524 14280 15552
rect 13009 15487 13067 15493
rect 13009 15453 13021 15487
rect 13055 15484 13067 15487
rect 13188 15484 13216 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 13055 15456 13216 15484
rect 13265 15487 13323 15493
rect 13055 15453 13067 15456
rect 13009 15447 13067 15453
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 13446 15484 13452 15496
rect 13311 15456 13452 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 17862 15484 17868 15496
rect 15703 15456 17868 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 17862 15444 17868 15456
rect 17920 15484 17926 15496
rect 18877 15487 18935 15493
rect 18877 15484 18889 15487
rect 17920 15456 18889 15484
rect 17920 15444 17926 15456
rect 18877 15453 18889 15456
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 13170 15376 13176 15428
rect 13228 15416 13234 15428
rect 15902 15419 15960 15425
rect 15902 15416 15914 15419
rect 13228 15388 15914 15416
rect 13228 15376 13234 15388
rect 15902 15385 15914 15388
rect 15948 15385 15960 15419
rect 18138 15416 18144 15428
rect 15902 15379 15960 15385
rect 17052 15388 18144 15416
rect 11882 15348 11888 15360
rect 11843 15320 11888 15348
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 17052 15357 17080 15388
rect 18138 15376 18144 15388
rect 18196 15376 18202 15428
rect 18632 15419 18690 15425
rect 18632 15385 18644 15419
rect 18678 15416 18690 15419
rect 19518 15416 19524 15428
rect 18678 15388 19524 15416
rect 18678 15385 18690 15388
rect 18632 15379 18690 15385
rect 19518 15376 19524 15388
rect 19576 15376 19582 15428
rect 13541 15351 13599 15357
rect 13541 15348 13553 15351
rect 13504 15320 13553 15348
rect 13504 15308 13510 15320
rect 13541 15317 13553 15320
rect 13587 15317 13599 15351
rect 13541 15311 13599 15317
rect 17037 15351 17095 15357
rect 17037 15317 17049 15351
rect 17083 15317 17095 15351
rect 17037 15311 17095 15317
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 17678 15348 17684 15360
rect 17543 15320 17684 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 5166 15104 5172 15156
rect 5224 15144 5230 15156
rect 5261 15147 5319 15153
rect 5261 15144 5273 15147
rect 5224 15116 5273 15144
rect 5224 15104 5230 15116
rect 5261 15113 5273 15116
rect 5307 15113 5319 15147
rect 5261 15107 5319 15113
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 6822 15144 6828 15156
rect 5767 15116 6828 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15144 7067 15147
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7055 15116 8033 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 8021 15113 8033 15116
rect 8067 15144 8079 15147
rect 8110 15144 8116 15156
rect 8067 15116 8116 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 16546 15116 16773 15144
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 9493 15079 9551 15085
rect 9493 15076 9505 15079
rect 7156 15048 9505 15076
rect 7156 15036 7162 15048
rect 9493 15045 9505 15048
rect 9539 15076 9551 15079
rect 9950 15076 9956 15088
rect 9539 15048 9956 15076
rect 9539 15045 9551 15048
rect 9493 15039 9551 15045
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 15964 15079 16022 15085
rect 15964 15045 15976 15079
rect 16010 15076 16022 15079
rect 16390 15076 16396 15088
rect 16010 15048 16396 15076
rect 16010 15045 16022 15048
rect 15964 15039 16022 15045
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 5626 15008 5632 15020
rect 5587 14980 5632 15008
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7650 15008 7656 15020
rect 6963 14980 7656 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 16206 15008 16212 15020
rect 16119 14980 16212 15008
rect 16206 14968 16212 14980
rect 16264 15008 16270 15020
rect 16546 15008 16574 15116
rect 16761 15113 16773 15116
rect 16807 15144 16819 15147
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 16807 15116 17233 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 17221 15113 17233 15116
rect 17267 15144 17279 15147
rect 17862 15144 17868 15156
rect 17267 15116 17868 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 20910 15079 20968 15085
rect 20910 15076 20922 15079
rect 20772 15048 20922 15076
rect 20772 15036 20778 15048
rect 20910 15045 20922 15048
rect 20956 15045 20968 15079
rect 20910 15039 20968 15045
rect 16264 14980 16574 15008
rect 21177 15011 21235 15017
rect 16264 14968 16270 14980
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 21266 15008 21272 15020
rect 21223 14980 21272 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 5905 14943 5963 14949
rect 5905 14909 5917 14943
rect 5951 14909 5963 14943
rect 5905 14903 5963 14909
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 14366 14940 14372 14952
rect 7239 14912 14372 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 5920 14872 5948 14903
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15194 14872 15200 14884
rect 5920 14844 15200 14872
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 4580 14776 6561 14804
rect 4580 14764 4586 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 7650 14804 7656 14816
rect 7611 14776 7656 14804
rect 6549 14767 6607 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 12986 14804 12992 14816
rect 9732 14776 12992 14804
rect 9732 14764 9738 14776
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14332 14776 14841 14804
rect 14332 14764 14338 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19576 14776 19809 14804
rect 19576 14764 19582 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 9784 14572 11621 14600
rect 9674 14532 9680 14544
rect 8036 14504 9680 14532
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 8036 14473 8064 14504
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 5684 14436 5733 14464
rect 5684 14424 5690 14436
rect 5721 14433 5733 14436
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 9784 14473 9812 14572
rect 11609 14569 11621 14572
rect 11655 14600 11667 14603
rect 11698 14600 11704 14612
rect 11655 14572 11704 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 16206 14600 16212 14612
rect 15887 14572 16212 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 9769 14467 9827 14473
rect 8260 14436 9628 14464
rect 8260 14424 8266 14436
rect 8205 14331 8263 14337
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8251 14300 8953 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 8110 14260 8116 14272
rect 8071 14232 8116 14260
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8573 14263 8631 14269
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 9490 14260 9496 14272
rect 8619 14232 9496 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9600 14260 9628 14436
rect 9769 14433 9781 14467
rect 9815 14433 9827 14467
rect 15473 14467 15531 14473
rect 9769 14427 9827 14433
rect 12912 14436 13492 14464
rect 9950 14396 9956 14408
rect 9911 14368 9956 14396
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14396 10103 14399
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10091 14368 10701 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 10060 14260 10088 14359
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12912 14396 12940 14436
rect 12492 14368 12940 14396
rect 12989 14399 13047 14405
rect 12492 14356 12498 14368
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 13464 14396 13492 14436
rect 15473 14433 15485 14467
rect 15519 14464 15531 14467
rect 15856 14464 15884 14563
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 19242 14600 19248 14612
rect 16316 14572 19248 14600
rect 15519 14436 15884 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 16316 14396 16344 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 21085 14603 21143 14609
rect 21085 14600 21097 14603
rect 19352 14572 21097 14600
rect 16390 14492 16396 14544
rect 16448 14532 16454 14544
rect 17497 14535 17555 14541
rect 17497 14532 17509 14535
rect 16448 14504 17509 14532
rect 16448 14492 16454 14504
rect 17497 14501 17509 14504
rect 17543 14501 17555 14535
rect 17497 14495 17555 14501
rect 19352 14473 19380 14572
rect 21085 14569 21097 14572
rect 21131 14600 21143 14603
rect 21266 14600 21272 14612
rect 21131 14572 21272 14600
rect 21131 14569 21143 14572
rect 21085 14563 21143 14569
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 18877 14467 18935 14473
rect 18877 14433 18889 14467
rect 18923 14464 18935 14467
rect 19337 14467 19395 14473
rect 19337 14464 19349 14467
rect 18923 14436 19349 14464
rect 18923 14433 18935 14436
rect 18877 14427 18935 14433
rect 19337 14433 19349 14436
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 13035 14368 13400 14396
rect 13464 14368 16344 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 12744 14331 12802 14337
rect 12744 14297 12756 14331
rect 12790 14328 12802 14331
rect 13078 14328 13084 14340
rect 12790 14300 13084 14328
rect 12790 14297 12802 14300
rect 12744 14291 12802 14297
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 9600 14232 10088 14260
rect 10413 14263 10471 14269
rect 10413 14229 10425 14263
rect 10459 14260 10471 14263
rect 10502 14260 10508 14272
rect 10459 14232 10508 14260
rect 10459 14229 10471 14232
rect 10413 14223 10471 14229
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 13372 14269 13400 14368
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 19593 14399 19651 14405
rect 19593 14396 19605 14399
rect 17368 14368 19605 14396
rect 17368 14356 17374 14368
rect 19593 14365 19605 14368
rect 19639 14396 19651 14399
rect 19978 14396 19984 14408
rect 19639 14368 19984 14396
rect 19639 14365 19651 14368
rect 19593 14359 19651 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 15194 14288 15200 14340
rect 15252 14337 15258 14340
rect 15252 14328 15264 14337
rect 15252 14300 15297 14328
rect 15252 14291 15264 14300
rect 15252 14288 15258 14291
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 17221 14331 17279 14337
rect 17221 14328 17233 14331
rect 15528 14300 17233 14328
rect 15528 14288 15534 14300
rect 17221 14297 17233 14300
rect 17267 14328 17279 14331
rect 18610 14331 18668 14337
rect 18610 14328 18622 14331
rect 17267 14300 18622 14328
rect 17267 14297 17279 14300
rect 17221 14291 17279 14297
rect 18610 14297 18622 14300
rect 18656 14297 18668 14331
rect 18610 14291 18668 14297
rect 13357 14263 13415 14269
rect 13357 14229 13369 14263
rect 13403 14260 13415 14263
rect 13446 14260 13452 14272
rect 13403 14232 13452 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13780 14232 14105 14260
rect 13780 14220 13786 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 20714 14260 20720 14272
rect 20675 14232 20720 14260
rect 14093 14223 14151 14229
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 4304 14028 6914 14056
rect 4304 14016 4310 14028
rect 6886 13920 6914 14028
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 8168 14028 8217 14056
rect 8168 14016 8174 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8205 14019 8263 14025
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 9306 14056 9312 14068
rect 9171 14028 9312 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 9456 14028 9597 14056
rect 9456 14016 9462 14028
rect 9585 14025 9597 14028
rect 9631 14056 9643 14059
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 9631 14028 10517 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 10744 14028 13553 14056
rect 10744 14016 10750 14028
rect 13541 14025 13553 14028
rect 13587 14056 13599 14059
rect 15470 14056 15476 14068
rect 13587 14028 15476 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 19061 14059 19119 14065
rect 19061 14025 19073 14059
rect 19107 14056 19119 14059
rect 20806 14056 20812 14068
rect 19107 14028 20812 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 20806 14016 20812 14028
rect 20864 14056 20870 14068
rect 21266 14056 21272 14068
rect 20864 14028 21272 14056
rect 20864 14016 20870 14028
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 7837 13991 7895 13997
rect 7837 13957 7849 13991
rect 7883 13988 7895 13991
rect 8573 13991 8631 13997
rect 8573 13988 8585 13991
rect 7883 13960 8585 13988
rect 7883 13957 7895 13960
rect 7837 13951 7895 13957
rect 8573 13957 8585 13960
rect 8619 13988 8631 13991
rect 9493 13991 9551 13997
rect 9493 13988 9505 13991
rect 8619 13960 9505 13988
rect 8619 13957 8631 13960
rect 8573 13951 8631 13957
rect 9493 13957 9505 13960
rect 9539 13988 9551 13991
rect 13446 13988 13452 14000
rect 9539 13960 10088 13988
rect 9539 13957 9551 13960
rect 9493 13951 9551 13957
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6886 13892 7205 13920
rect 7193 13889 7205 13892
rect 7239 13920 7251 13923
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7239 13892 7757 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 9600 13892 9812 13920
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13821 7711 13855
rect 9600 13852 9628 13892
rect 7653 13815 7711 13821
rect 9508 13824 9628 13852
rect 9677 13855 9735 13861
rect 7668 13784 7696 13815
rect 9508 13784 9536 13824
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9692 13784 9720 13815
rect 7668 13756 9536 13784
rect 9600 13756 9720 13784
rect 9784 13784 9812 13892
rect 10060 13864 10088 13960
rect 12176 13960 13452 13988
rect 12176 13929 12204 13960
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12417 13923 12475 13929
rect 12417 13920 12429 13923
rect 12161 13883 12219 13889
rect 12268 13892 12429 13920
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 10100 13824 10149 13852
rect 10100 13812 10106 13824
rect 10137 13821 10149 13824
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12268 13852 12296 13892
rect 12417 13889 12429 13892
rect 12463 13889 12475 13923
rect 12417 13883 12475 13889
rect 11756 13824 12296 13852
rect 11756 13812 11762 13824
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13504 13824 13921 13852
rect 13504 13812 13510 13824
rect 13909 13821 13921 13824
rect 13955 13852 13967 13855
rect 16206 13852 16212 13864
rect 13955 13824 16212 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 20070 13852 20076 13864
rect 19392 13824 20076 13852
rect 19392 13812 19398 13824
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 11882 13784 11888 13796
rect 9784 13756 11888 13784
rect 9600 13728 9628 13756
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 16390 13784 16396 13796
rect 13464 13756 16396 13784
rect 9582 13676 9588 13728
rect 9640 13676 9646 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 13464 13716 13492 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 11664 13688 13492 13716
rect 11664 13676 11670 13688
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 19702 13716 19708 13728
rect 17644 13688 19708 13716
rect 17644 13676 17650 13688
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 21174 13676 21180 13728
rect 21232 13716 21238 13728
rect 21269 13719 21327 13725
rect 21269 13716 21281 13719
rect 21232 13688 21281 13716
rect 21232 13676 21238 13688
rect 21269 13685 21281 13688
rect 21315 13685 21327 13719
rect 21269 13679 21327 13685
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 4488 13484 5917 13512
rect 4488 13472 4494 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 5905 13475 5963 13481
rect 5920 13308 5948 13475
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 7340 13484 7389 13512
rect 7340 13472 7346 13484
rect 7377 13481 7389 13484
rect 7423 13512 7435 13515
rect 7742 13512 7748 13524
rect 7423 13484 7748 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 7742 13472 7748 13484
rect 7800 13512 7806 13524
rect 8018 13512 8024 13524
rect 7800 13484 8024 13512
rect 7800 13472 7806 13484
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 9766 13512 9772 13524
rect 9723 13484 9772 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 13446 13512 13452 13524
rect 11716 13484 12664 13512
rect 13407 13484 13452 13512
rect 11606 13444 11612 13456
rect 6886 13416 11612 13444
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6886 13376 6914 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 6503 13348 6914 13376
rect 9125 13379 9183 13385
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 9125 13345 9137 13379
rect 9171 13376 9183 13379
rect 11716 13376 11744 13484
rect 12636 13444 12664 13484
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 16264 13484 16405 13512
rect 16264 13472 16270 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 16393 13475 16451 13481
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 18104 13484 21005 13512
rect 18104 13472 18110 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 12636 13416 13584 13444
rect 9171 13348 11744 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 5920 13280 6561 13308
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13308 6699 13311
rect 7282 13308 7288 13320
rect 6687 13280 7288 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 10870 13308 10876 13320
rect 9263 13280 10876 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13308 11759 13311
rect 13446 13308 13452 13320
rect 11747 13280 13452 13308
rect 11747 13277 11759 13280
rect 11701 13271 11759 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13556 13308 13584 13416
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13376 16175 13379
rect 16224 13376 16252 13472
rect 16163 13348 16252 13376
rect 20625 13379 20683 13385
rect 16163 13345 16175 13348
rect 16117 13339 16175 13345
rect 20625 13345 20637 13379
rect 20671 13376 20683 13379
rect 20806 13376 20812 13388
rect 20671 13348 20812 13376
rect 20671 13345 20683 13348
rect 20625 13339 20683 13345
rect 17586 13308 17592 13320
rect 13556 13280 17592 13308
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 17966 13311 18024 13317
rect 17966 13277 17978 13311
rect 18012 13277 18024 13311
rect 17966 13271 18024 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18414 13308 18420 13320
rect 18279 13280 18420 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 8294 13240 8300 13252
rect 6788 13212 8300 13240
rect 6788 13200 6794 13212
rect 8294 13200 8300 13212
rect 8352 13240 8358 13252
rect 9309 13243 9367 13249
rect 9309 13240 9321 13243
rect 8352 13212 9321 13240
rect 8352 13200 8358 13212
rect 9309 13209 9321 13212
rect 9355 13240 9367 13243
rect 9953 13243 10011 13249
rect 9953 13240 9965 13243
rect 9355 13212 9965 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 9953 13209 9965 13212
rect 9999 13209 10011 13243
rect 9953 13203 10011 13209
rect 11968 13243 12026 13249
rect 11968 13209 11980 13243
rect 12014 13240 12026 13243
rect 12434 13240 12440 13252
rect 12014 13212 12440 13240
rect 12014 13209 12026 13212
rect 11968 13203 12026 13209
rect 12434 13200 12440 13212
rect 12492 13240 12498 13252
rect 13722 13240 13728 13252
rect 12492 13212 13728 13240
rect 12492 13200 12498 13212
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 15850 13243 15908 13249
rect 15850 13240 15862 13243
rect 15620 13212 15862 13240
rect 15620 13200 15626 13212
rect 15850 13209 15862 13212
rect 15896 13209 15908 13243
rect 17972 13240 18000 13271
rect 18414 13268 18420 13280
rect 18472 13308 18478 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 18472 13280 18613 13308
rect 18472 13268 18478 13280
rect 18601 13277 18613 13280
rect 18647 13308 18659 13311
rect 20640 13308 20668 13339
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 21174 13308 21180 13320
rect 18647 13280 20668 13308
rect 21135 13280 21180 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 18046 13240 18052 13252
rect 15850 13203 15908 13209
rect 15948 13212 17908 13240
rect 17972 13212 18052 13240
rect 7006 13172 7012 13184
rect 6967 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 10410 13172 10416 13184
rect 10371 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 13078 13172 13084 13184
rect 12991 13144 13084 13172
rect 13078 13132 13084 13144
rect 13136 13172 13142 13184
rect 13354 13172 13360 13184
rect 13136 13144 13360 13172
rect 13136 13132 13142 13144
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13538 13132 13544 13184
rect 13596 13172 13602 13184
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 13596 13144 14749 13172
rect 13596 13132 13602 13144
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 14737 13135 14795 13141
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15948 13172 15976 13212
rect 14884 13144 15976 13172
rect 14884 13132 14890 13144
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16080 13144 16865 13172
rect 16080 13132 16086 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 17880 13172 17908 13212
rect 18046 13200 18052 13212
rect 18104 13200 18110 13252
rect 20358 13243 20416 13249
rect 20358 13240 20370 13243
rect 19812 13212 20370 13240
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 17880 13144 19257 13172
rect 16853 13135 16911 13141
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19812 13172 19840 13212
rect 20358 13209 20370 13212
rect 20404 13209 20416 13243
rect 20358 13203 20416 13209
rect 19392 13144 19840 13172
rect 19392 13132 19398 13144
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 7616 12940 10057 12968
rect 7616 12928 7622 12940
rect 10045 12937 10057 12940
rect 10091 12937 10103 12971
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 10045 12931 10103 12937
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 13446 12968 13452 12980
rect 10560 12940 10605 12968
rect 13407 12940 13452 12968
rect 10560 12928 10566 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 18414 12968 18420 12980
rect 18375 12940 18420 12968
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 12814 12903 12872 12909
rect 12814 12900 12826 12903
rect 11204 12872 12826 12900
rect 11204 12860 11210 12872
rect 12814 12869 12826 12872
rect 12860 12869 12872 12903
rect 12814 12863 12872 12869
rect 12526 12832 12532 12844
rect 10704 12804 12532 12832
rect 10704 12773 10732 12804
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13464 12832 13492 12928
rect 18432 12900 18460 12928
rect 16684 12872 18460 12900
rect 16684 12841 16712 12872
rect 20806 12860 20812 12912
rect 20864 12900 20870 12912
rect 21266 12900 21272 12912
rect 20864 12872 21272 12900
rect 20864 12860 20870 12872
rect 21266 12860 21272 12872
rect 21324 12900 21330 12912
rect 21324 12872 21404 12900
rect 21324 12860 21330 12872
rect 21376 12841 21404 12872
rect 13127 12804 13492 12832
rect 16669 12835 16727 12841
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 16669 12801 16681 12835
rect 16715 12801 16727 12835
rect 16925 12835 16983 12841
rect 16925 12832 16937 12835
rect 16669 12795 16727 12801
rect 16776 12804 16937 12832
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12733 10747 12767
rect 10689 12727 10747 12733
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 16776 12764 16804 12804
rect 16925 12801 16937 12804
rect 16971 12801 16983 12835
rect 21094 12835 21152 12841
rect 21094 12832 21106 12835
rect 16925 12795 16983 12801
rect 19628 12804 21106 12832
rect 15528 12736 16804 12764
rect 15528 12724 15534 12736
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 19628 12705 19656 12804
rect 21094 12801 21106 12804
rect 21140 12801 21152 12835
rect 21094 12795 21152 12801
rect 21361 12835 21419 12841
rect 21361 12801 21373 12835
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 19613 12699 19671 12705
rect 19613 12696 19625 12699
rect 17736 12668 19625 12696
rect 17736 12656 17742 12668
rect 19613 12665 19625 12668
rect 19659 12665 19671 12699
rect 19613 12659 19671 12665
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 9640 12600 11713 12628
rect 9640 12588 9646 12600
rect 11701 12597 11713 12600
rect 11747 12628 11759 12631
rect 13814 12628 13820 12640
rect 11747 12600 13820 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 17954 12628 17960 12640
rect 15712 12600 17960 12628
rect 15712 12588 15718 12600
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 18874 12628 18880 12640
rect 18095 12600 18880 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 18874 12588 18880 12600
rect 18932 12628 18938 12640
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 18932 12600 19073 12628
rect 18932 12588 18938 12600
rect 19061 12597 19073 12600
rect 19107 12628 19119 12631
rect 19242 12628 19248 12640
rect 19107 12600 19248 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19978 12628 19984 12640
rect 19939 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 16022 12424 16028 12436
rect 12400 12396 16028 12424
rect 12400 12384 12406 12396
rect 16022 12384 16028 12396
rect 16080 12384 16086 12436
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 11238 12288 11244 12300
rect 10091 12260 11244 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10192 12192 10241 12220
rect 10192 12180 10198 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 17218 12220 17224 12232
rect 17000 12192 17224 12220
rect 17000 12180 17006 12192
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 19978 12220 19984 12232
rect 18472 12192 19984 12220
rect 18472 12180 18478 12192
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 21266 12220 21272 12232
rect 21227 12192 21272 12220
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 15194 12152 15200 12164
rect 12768 12124 15200 12152
rect 12768 12112 12774 12124
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 15286 12112 15292 12164
rect 15344 12152 15350 12164
rect 21002 12155 21060 12161
rect 21002 12152 21014 12155
rect 15344 12124 21014 12152
rect 15344 12112 15350 12124
rect 21002 12121 21014 12124
rect 21048 12121 21060 12155
rect 21002 12115 21060 12121
rect 5997 12087 6055 12093
rect 5997 12053 6009 12087
rect 6043 12084 6055 12087
rect 6730 12084 6736 12096
rect 6043 12056 6736 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 14274 12084 14280 12096
rect 6880 12056 14280 12084
rect 6880 12044 6886 12056
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 18414 12084 18420 12096
rect 16080 12056 18420 12084
rect 16080 12044 16086 12056
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18690 12044 18696 12096
rect 18748 12084 18754 12096
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 18748 12056 19533 12084
rect 18748 12044 18754 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 19889 12087 19947 12093
rect 19889 12084 19901 12087
rect 19852 12056 19901 12084
rect 19852 12044 19858 12056
rect 19889 12053 19901 12056
rect 19935 12053 19947 12087
rect 19889 12047 19947 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 6730 11880 6736 11892
rect 6691 11852 6736 11880
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7147 11852 12434 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 6641 11815 6699 11821
rect 6641 11781 6653 11815
rect 6687 11812 6699 11815
rect 7006 11812 7012 11824
rect 6687 11784 7012 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 12406 11812 12434 11852
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 17034 11880 17040 11892
rect 12860 11852 17040 11880
rect 12860 11840 12866 11852
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 17144 11852 18981 11880
rect 14550 11812 14556 11824
rect 12406 11784 14556 11812
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 17144 11812 17172 11852
rect 18969 11849 18981 11852
rect 19015 11880 19027 11883
rect 19058 11880 19064 11892
rect 19015 11852 19064 11880
rect 19015 11849 19027 11852
rect 18969 11843 19027 11849
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 15252 11784 17172 11812
rect 15252 11772 15258 11784
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 17920 11784 18644 11812
rect 17920 11772 17926 11784
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 14113 11747 14171 11753
rect 14113 11744 14125 11747
rect 13688 11716 14125 11744
rect 13688 11704 13694 11716
rect 14113 11713 14125 11716
rect 14159 11713 14171 11747
rect 14113 11707 14171 11713
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 14415 11716 14780 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 6549 11679 6607 11685
rect 6549 11645 6561 11679
rect 6595 11676 6607 11679
rect 6822 11676 6828 11688
rect 6595 11648 6828 11676
rect 6595 11645 6607 11648
rect 6549 11639 6607 11645
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 11146 11568 11152 11620
rect 11204 11608 11210 11620
rect 13354 11608 13360 11620
rect 11204 11580 13360 11608
rect 11204 11568 11210 11580
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 12802 11540 12808 11552
rect 7340 11512 12808 11540
rect 7340 11500 7346 11512
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 12986 11540 12992 11552
rect 12947 11512 12992 11540
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 14752 11549 14780 11716
rect 18414 11704 18420 11756
rect 18472 11753 18478 11756
rect 18472 11744 18484 11753
rect 18616 11744 18644 11784
rect 18690 11772 18696 11824
rect 18748 11812 18754 11824
rect 18748 11784 20392 11812
rect 18748 11772 18754 11784
rect 19794 11744 19800 11756
rect 18472 11716 18517 11744
rect 18616 11716 19800 11744
rect 18472 11707 18484 11716
rect 18472 11704 18478 11707
rect 19794 11704 19800 11716
rect 19852 11744 19858 11756
rect 20364 11753 20392 11784
rect 20082 11747 20140 11753
rect 20082 11744 20094 11747
rect 19852 11716 20094 11744
rect 19852 11704 19858 11716
rect 20082 11713 20094 11716
rect 20128 11713 20140 11747
rect 20082 11707 20140 11713
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11744 20407 11747
rect 20625 11747 20683 11753
rect 20625 11744 20637 11747
rect 20395 11716 20637 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 20625 11713 20637 11716
rect 20671 11744 20683 11747
rect 20898 11744 20904 11756
rect 20671 11716 20904 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 20898 11704 20904 11716
rect 20956 11744 20962 11756
rect 21266 11744 21272 11756
rect 20956 11716 21272 11744
rect 20956 11704 20962 11716
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 18690 11676 18696 11688
rect 18651 11648 18696 11676
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15010 11540 15016 11552
rect 14783 11512 15016 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 17402 11540 17408 11552
rect 17359 11512 17408 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 12894 11336 12900 11348
rect 10980 11308 12900 11336
rect 9585 11203 9643 11209
rect 9585 11169 9597 11203
rect 9631 11200 9643 11203
rect 10980 11200 11008 11308
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 13412 11308 15945 11336
rect 13412 11296 13418 11308
rect 15933 11305 15945 11308
rect 15979 11305 15991 11339
rect 15933 11299 15991 11305
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 20530 11336 20536 11348
rect 17736 11308 20536 11336
rect 17736 11296 17742 11308
rect 20530 11296 20536 11308
rect 20588 11336 20594 11348
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 20588 11308 20637 11336
rect 20588 11296 20594 11308
rect 20625 11305 20637 11308
rect 20671 11305 20683 11339
rect 20898 11336 20904 11348
rect 20859 11308 20904 11336
rect 20625 11299 20683 11305
rect 20898 11296 20904 11308
rect 20956 11296 20962 11348
rect 15470 11268 15476 11280
rect 15431 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 9631 11172 11008 11200
rect 9631 11169 9643 11172
rect 9585 11163 9643 11169
rect 19058 11160 19064 11212
rect 19116 11200 19122 11212
rect 19116 11172 19380 11200
rect 19116 11160 19122 11172
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 12713 11135 12771 11141
rect 9723 11104 12664 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 9769 11067 9827 11073
rect 9769 11033 9781 11067
rect 9815 11064 9827 11067
rect 10413 11067 10471 11073
rect 10413 11064 10425 11067
rect 9815 11036 10425 11064
rect 9815 11033 9827 11036
rect 9769 11027 9827 11033
rect 10413 11033 10425 11036
rect 10459 11033 10471 11067
rect 10413 11027 10471 11033
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 12342 11064 12348 11076
rect 11848 11036 12348 11064
rect 11848 11024 11854 11036
rect 12342 11024 12348 11036
rect 12400 11064 12406 11076
rect 12446 11067 12504 11073
rect 12446 11064 12458 11067
rect 12400 11036 12458 11064
rect 12400 11024 12406 11036
rect 12446 11033 12458 11036
rect 12492 11033 12504 11067
rect 12636 11064 12664 11104
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12759 11104 13093 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 13081 11101 13093 11104
rect 13127 11132 13139 11135
rect 13262 11132 13268 11144
rect 13127 11104 13268 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13262 11092 13268 11104
rect 13320 11132 13326 11144
rect 13446 11132 13452 11144
rect 13320 11104 13452 11132
rect 13320 11092 13326 11104
rect 13446 11092 13452 11104
rect 13504 11132 13510 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13504 11104 14105 11132
rect 13504 11092 13510 11104
rect 14093 11101 14105 11104
rect 14139 11132 14151 11135
rect 14139 11104 15056 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 15028 11076 15056 11104
rect 17034 11092 17040 11144
rect 17092 11141 17098 11144
rect 17092 11132 17104 11141
rect 17310 11132 17316 11144
rect 17092 11104 17172 11132
rect 17271 11104 17316 11132
rect 17092 11095 17104 11104
rect 17092 11092 17098 11095
rect 12636 11036 13768 11064
rect 12446 11027 12504 11033
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11333 10999 11391 11005
rect 11333 10996 11345 10999
rect 11112 10968 11345 10996
rect 11112 10956 11118 10968
rect 11333 10965 11345 10968
rect 11379 10965 11391 10999
rect 11333 10959 11391 10965
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13538 10996 13544 11008
rect 12952 10968 13544 10996
rect 12952 10956 12958 10968
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 13740 10996 13768 11036
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14338 11067 14396 11073
rect 14338 11064 14350 11067
rect 13872 11036 14350 11064
rect 13872 11024 13878 11036
rect 14338 11033 14350 11036
rect 14384 11033 14396 11067
rect 14338 11027 14396 11033
rect 15010 11024 15016 11076
rect 15068 11024 15074 11076
rect 17144 11064 17172 11104
rect 17310 11092 17316 11104
rect 17368 11132 17374 11144
rect 17589 11135 17647 11141
rect 17589 11132 17601 11135
rect 17368 11104 17601 11132
rect 17368 11092 17374 11104
rect 17589 11101 17601 11104
rect 17635 11132 17647 11135
rect 18690 11132 18696 11144
rect 17635 11104 18696 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 18690 11092 18696 11104
rect 18748 11132 18754 11144
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 18748 11104 18797 11132
rect 18748 11092 18754 11104
rect 18785 11101 18797 11104
rect 18831 11132 18843 11135
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18831 11104 19257 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19352 11132 19380 11172
rect 19501 11135 19559 11141
rect 19501 11132 19513 11135
rect 19352 11104 19513 11132
rect 19245 11095 19303 11101
rect 19501 11101 19513 11104
rect 19547 11101 19559 11135
rect 19501 11095 19559 11101
rect 19150 11064 19156 11076
rect 17144 11036 19156 11064
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 15194 10996 15200 11008
rect 13740 10968 15200 10996
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 6871 10764 7573 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 7561 10755 7619 10761
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8202 10792 8208 10804
rect 7975 10764 8208 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 12894 10792 12900 10804
rect 8772 10764 12900 10792
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 8021 10727 8079 10733
rect 8021 10724 8033 10727
rect 7432 10696 8033 10724
rect 7432 10684 7438 10696
rect 8021 10693 8033 10696
rect 8067 10693 8079 10727
rect 8021 10687 8079 10693
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7098 10656 7104 10668
rect 6963 10628 7104 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 8772 10656 8800 10764
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13262 10792 13268 10804
rect 13223 10764 13268 10792
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 15657 10795 15715 10801
rect 15657 10761 15669 10795
rect 15703 10792 15715 10795
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15703 10764 15945 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 13280 10724 13308 10752
rect 11532 10696 13308 10724
rect 11532 10665 11560 10696
rect 8128 10628 8800 10656
rect 11517 10659 11575 10665
rect 6733 10591 6791 10597
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 8128 10588 8156 10628
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11773 10659 11831 10665
rect 11773 10656 11785 10659
rect 11517 10619 11575 10625
rect 11624 10628 11785 10656
rect 6779 10560 8156 10588
rect 8205 10591 8263 10597
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 9309 10591 9367 10597
rect 8251 10560 9260 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 8110 10452 8116 10464
rect 7331 10424 8116 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8573 10455 8631 10461
rect 8573 10452 8585 10455
rect 8260 10424 8585 10452
rect 8260 10412 8266 10424
rect 8573 10421 8585 10424
rect 8619 10421 8631 10455
rect 9232 10452 9260 10560
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 9398 10588 9404 10600
rect 9355 10560 9404 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11624 10588 11652 10628
rect 11773 10625 11785 10628
rect 11819 10625 11831 10659
rect 11773 10619 11831 10625
rect 14734 10616 14740 10668
rect 14792 10665 14798 10668
rect 14792 10656 14804 10665
rect 14792 10628 14837 10656
rect 14792 10619 14804 10628
rect 14792 10616 14798 10619
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 15672 10656 15700 10755
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 17460 10764 18644 10792
rect 17460 10752 17466 10764
rect 17310 10684 17316 10736
rect 17368 10724 17374 10736
rect 18509 10727 18567 10733
rect 18509 10724 18521 10727
rect 17368 10696 18521 10724
rect 17368 10684 17374 10696
rect 15068 10628 15700 10656
rect 15068 10616 15074 10628
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 18248 10665 18276 10696
rect 18509 10693 18521 10696
rect 18555 10693 18567 10727
rect 18509 10687 18567 10693
rect 17966 10659 18024 10665
rect 17966 10656 17978 10659
rect 16908 10628 17978 10656
rect 16908 10616 16914 10628
rect 17966 10625 17978 10628
rect 18012 10625 18024 10659
rect 17966 10619 18024 10625
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10625 18291 10659
rect 18616 10656 18644 10764
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19208 10764 19809 10792
rect 19208 10752 19214 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 20916 10724 20944 10752
rect 20916 10696 21220 10724
rect 21192 10665 21220 10696
rect 20910 10659 20968 10665
rect 20910 10656 20922 10659
rect 18616 10628 20922 10656
rect 18233 10619 18291 10625
rect 20910 10625 20922 10628
rect 20956 10625 20968 10659
rect 20910 10619 20968 10625
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 21266 10656 21272 10668
rect 21223 10628 21272 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 11112 10560 11652 10588
rect 11112 10548 11118 10560
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10520 12955 10523
rect 12943 10492 13768 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 12912 10452 12940 10483
rect 13630 10452 13636 10464
rect 9232 10424 12940 10452
rect 13591 10424 13636 10452
rect 8573 10415 8631 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 13740 10452 13768 10492
rect 15562 10452 15568 10464
rect 13740 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16482 10412 16488 10464
rect 16540 10452 16546 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16540 10424 16865 10452
rect 16540 10412 16546 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 12710 10248 12716 10260
rect 9232 10220 12716 10248
rect 7098 10112 7104 10124
rect 7059 10084 7104 10112
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 9232 10121 9260 10220
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 15197 10251 15255 10257
rect 15197 10217 15209 10251
rect 15243 10248 15255 10251
rect 15286 10248 15292 10260
rect 15243 10220 15292 10248
rect 15243 10217 15255 10220
rect 15197 10211 15255 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 10413 10115 10471 10121
rect 9217 10075 9275 10081
rect 9692 10084 10364 10112
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 9398 10044 9404 10056
rect 9359 10016 9404 10044
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 8389 9979 8447 9985
rect 8389 9945 8401 9979
rect 8435 9976 8447 9979
rect 9692 9976 9720 10084
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 8435 9948 9720 9976
rect 9784 10016 10149 10044
rect 8435 9945 8447 9948
rect 8389 9939 8447 9945
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9784 9917 9812 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10336 10044 10364 10084
rect 10413 10081 10425 10115
rect 10459 10112 10471 10115
rect 10594 10112 10600 10124
rect 10459 10084 10600 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 13280 10112 13308 10208
rect 13035 10084 13308 10112
rect 16577 10115 16635 10121
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 16623 10084 17233 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 17221 10081 17233 10084
rect 17267 10112 17279 10115
rect 17310 10112 17316 10124
rect 17267 10084 17316 10112
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 12250 10044 12256 10056
rect 10336 10016 12256 10044
rect 10137 10007 10195 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12733 10047 12791 10053
rect 12733 10013 12745 10047
rect 12779 10044 12791 10047
rect 12894 10044 12900 10056
rect 12779 10016 12900 10044
rect 12779 10013 12791 10016
rect 12733 10007 12791 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 16321 10047 16379 10053
rect 16321 10013 16333 10047
rect 16367 10044 16379 10047
rect 16482 10044 16488 10056
rect 16367 10016 16488 10044
rect 16367 10013 16379 10016
rect 16321 10007 16379 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9877 9827 9911
rect 9769 9871 9827 9877
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 11609 9911 11667 9917
rect 11609 9908 11621 9911
rect 11296 9880 11621 9908
rect 11296 9868 11302 9880
rect 11609 9877 11621 9880
rect 11655 9908 11667 9911
rect 11698 9908 11704 9920
rect 11655 9880 11704 9908
rect 11655 9877 11667 9880
rect 11609 9871 11667 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 16850 9908 16856 9920
rect 15068 9880 16856 9908
rect 15068 9868 15074 9880
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 17218 9704 17224 9716
rect 9364 9676 17224 9704
rect 9364 9664 9370 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 6696 9608 7389 9636
rect 6696 9596 6702 9608
rect 7377 9605 7389 9608
rect 7423 9636 7435 9639
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 7423 9608 8217 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 13872 9608 15516 9636
rect 13872 9596 13878 9608
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7708 9540 8125 9568
rect 7708 9528 7714 9540
rect 8113 9537 8125 9540
rect 8159 9568 8171 9571
rect 8662 9568 8668 9580
rect 8159 9540 8668 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8662 9528 8668 9540
rect 8720 9568 8726 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8720 9540 8769 9568
rect 8720 9528 8726 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 12250 9568 12256 9580
rect 12211 9540 12256 9568
rect 8757 9531 8815 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 15102 9528 15108 9580
rect 15160 9568 15166 9580
rect 15488 9577 15516 9608
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 15160 9540 15209 9568
rect 15160 9528 15166 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 20530 9568 20536 9580
rect 20491 9540 20536 9568
rect 19705 9531 19763 9537
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 8389 9503 8447 9509
rect 6604 9472 7880 9500
rect 6604 9460 6610 9472
rect 5718 9392 5724 9444
rect 5776 9432 5782 9444
rect 7745 9435 7803 9441
rect 7745 9432 7757 9435
rect 5776 9404 7757 9432
rect 5776 9392 5782 9404
rect 7745 9401 7757 9404
rect 7791 9401 7803 9435
rect 7852 9432 7880 9472
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 11238 9500 11244 9512
rect 8435 9472 11244 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9500 15071 9503
rect 19720 9500 19748 9531
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 21358 9568 21364 9580
rect 21319 9540 21364 9568
rect 21358 9528 21364 9540
rect 21416 9528 21422 9580
rect 15059 9472 19748 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 12342 9432 12348 9444
rect 7852 9404 12348 9432
rect 7745 9395 7803 9401
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 12437 9435 12495 9441
rect 12437 9401 12449 9435
rect 12483 9432 12495 9435
rect 14458 9432 14464 9444
rect 12483 9404 14464 9432
rect 12483 9401 12495 9404
rect 12437 9395 12495 9401
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 15654 9432 15660 9444
rect 15615 9404 15660 9432
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 19886 9432 19892 9444
rect 19847 9404 19892 9432
rect 19886 9392 19892 9404
rect 19944 9392 19950 9444
rect 20622 9392 20628 9444
rect 20680 9432 20686 9444
rect 20717 9435 20775 9441
rect 20717 9432 20729 9435
rect 20680 9404 20729 9432
rect 20680 9392 20686 9404
rect 20717 9401 20729 9404
rect 20763 9401 20775 9435
rect 20717 9395 20775 9401
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 17126 9364 17132 9376
rect 12768 9336 17132 9364
rect 12768 9324 12774 9336
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 21174 9364 21180 9376
rect 21135 9336 21180 9364
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 5552 9132 7021 9160
rect 5552 9033 5580 9132
rect 7009 9129 7021 9132
rect 7055 9160 7067 9163
rect 10686 9160 10692 9172
rect 7055 9132 10692 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 14182 9160 14188 9172
rect 12400 9132 14188 9160
rect 12400 9120 12406 9132
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14476 9132 15240 9160
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9061 6239 9095
rect 14476 9092 14504 9132
rect 6181 9055 6239 9061
rect 9232 9064 14504 9092
rect 15212 9092 15240 9132
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 17218 9160 17224 9172
rect 15344 9132 15389 9160
rect 17179 9132 17224 9160
rect 15344 9120 15350 9132
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 18322 9120 18328 9172
rect 18380 9160 18386 9172
rect 19429 9163 19487 9169
rect 19429 9160 19441 9163
rect 18380 9132 19441 9160
rect 18380 9120 18386 9132
rect 19429 9129 19441 9132
rect 19475 9129 19487 9163
rect 20438 9160 20444 9172
rect 20399 9132 20444 9160
rect 19429 9123 19487 9129
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 15212 9064 19288 9092
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 8993 5595 9027
rect 5718 9024 5724 9036
rect 5679 8996 5724 9024
rect 5537 8987 5595 8993
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 6196 8956 6224 9055
rect 9232 9033 9260 9064
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 10836 8996 13093 9024
rect 10836 8984 10842 8996
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16390 9024 16396 9036
rect 15979 8996 16396 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 17862 9024 17868 9036
rect 17823 8996 17868 9024
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 6196 8928 8953 8956
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13320 8928 13369 8956
rect 13320 8916 13326 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 14550 8956 14556 8968
rect 14511 8928 14556 8956
rect 13357 8919 13415 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15620 8928 15761 8956
rect 15620 8916 15626 8928
rect 15749 8925 15761 8928
rect 15795 8956 15807 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 15795 8928 16865 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 16942 8956 16948 8968
rect 16899 8928 16948 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 16942 8916 16948 8928
rect 17000 8956 17006 8968
rect 19260 8965 19288 9064
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 17000 8928 17693 8956
rect 17000 8916 17006 8928
rect 17681 8925 17693 8928
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 19245 8959 19303 8965
rect 19245 8925 19257 8959
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 21358 8956 21364 8968
rect 20671 8928 21036 8956
rect 21319 8928 21364 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 5813 8891 5871 8897
rect 5813 8857 5825 8891
rect 5859 8888 5871 8891
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 5859 8860 6469 8888
rect 5859 8857 5871 8860
rect 5813 8851 5871 8857
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 14829 8891 14887 8897
rect 11940 8860 14780 8888
rect 11940 8848 11946 8860
rect 12452 8829 12480 8860
rect 12437 8823 12495 8829
rect 12437 8789 12449 8823
rect 12483 8820 12495 8823
rect 14752 8820 14780 8860
rect 14829 8857 14841 8891
rect 14875 8888 14887 8891
rect 19812 8888 19840 8919
rect 14875 8860 19840 8888
rect 14875 8857 14887 8860
rect 14829 8851 14887 8857
rect 21008 8832 21036 8928
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 15562 8820 15568 8832
rect 12483 8792 12517 8820
rect 14752 8792 15568 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8820 15715 8823
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 15703 8792 16405 8820
rect 15703 8789 15715 8792
rect 15657 8783 15715 8789
rect 16393 8789 16405 8792
rect 16439 8820 16451 8823
rect 17494 8820 17500 8832
rect 16439 8792 17500 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 18322 8820 18328 8832
rect 17635 8792 18328 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19981 8823 20039 8829
rect 19981 8820 19993 8823
rect 19024 8792 19993 8820
rect 19024 8780 19030 8792
rect 19981 8789 19993 8792
rect 20027 8789 20039 8823
rect 20990 8820 20996 8832
rect 20951 8792 20996 8820
rect 19981 8783 20039 8789
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 5868 8588 6745 8616
rect 5868 8576 5874 8588
rect 6733 8585 6745 8588
rect 6779 8616 6791 8619
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 6779 8588 7389 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9263 8588 9873 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 9861 8579 9919 8585
rect 10704 8588 11805 8616
rect 10704 8560 10732 8588
rect 11793 8585 11805 8588
rect 11839 8616 11851 8619
rect 11882 8616 11888 8628
rect 11839 8588 11888 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 13262 8616 13268 8628
rect 12299 8588 12434 8616
rect 13223 8588 13268 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 10321 8551 10379 8557
rect 10321 8548 10333 8551
rect 7892 8520 10333 8548
rect 7892 8508 7898 8520
rect 10321 8517 10333 8520
rect 10367 8548 10379 8551
rect 10686 8548 10692 8560
rect 10367 8520 10692 8548
rect 10367 8517 10379 8520
rect 10321 8511 10379 8517
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 11146 8548 11152 8560
rect 11072 8520 11152 8548
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 9582 8480 9588 8492
rect 7515 8452 8156 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7282 8412 7288 8424
rect 7243 8384 7288 8412
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 8128 8356 8156 8452
rect 8956 8452 9588 8480
rect 8956 8421 8984 8452
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10275 8452 10885 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10873 8449 10885 8452
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 8941 8375 8999 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 10410 8372 10416 8424
rect 10468 8412 10474 8424
rect 11072 8412 11100 8520
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 12406 8548 12434 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 15102 8616 15108 8628
rect 15063 8588 15108 8616
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 17497 8619 17555 8625
rect 17497 8585 17509 8619
rect 17543 8616 17555 8619
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17543 8588 18061 8616
rect 17543 8585 17555 8588
rect 17497 8579 17555 8585
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 18049 8579 18107 8585
rect 18506 8576 18512 8628
rect 18564 8616 18570 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 18564 8588 19257 8616
rect 18564 8576 18570 8588
rect 19245 8585 19257 8588
rect 19291 8585 19303 8619
rect 19245 8579 19303 8585
rect 19889 8619 19947 8625
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 20070 8616 20076 8628
rect 19935 8588 20076 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 20438 8616 20444 8628
rect 20399 8588 20444 8616
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 14737 8551 14795 8557
rect 14737 8548 14749 8551
rect 12406 8520 14749 8548
rect 14737 8517 14749 8520
rect 14783 8517 14795 8551
rect 14737 8511 14795 8517
rect 15657 8551 15715 8557
rect 15657 8517 15669 8551
rect 15703 8548 15715 8551
rect 20714 8548 20720 8560
rect 15703 8520 19104 8548
rect 15703 8517 15715 8520
rect 15657 8511 15715 8517
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 12943 8452 13553 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 15930 8480 15936 8492
rect 15891 8452 15936 8480
rect 13541 8443 13599 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 18046 8480 18052 8492
rect 17451 8452 18052 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8480 18475 8483
rect 18874 8480 18880 8492
rect 18463 8452 18880 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19076 8489 19104 8520
rect 19628 8520 20720 8548
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 10468 8384 11100 8412
rect 10468 8372 10474 8384
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11204 8384 11621 8412
rect 11204 8372 11210 8384
rect 11609 8381 11621 8384
rect 11655 8412 11667 8415
rect 12710 8412 12716 8424
rect 11655 8384 12434 8412
rect 12671 8384 12716 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 8110 8344 8116 8356
rect 8071 8316 8116 8344
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 12406 8344 12434 8384
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 14366 8412 14372 8424
rect 12851 8384 14372 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14461 8415 14519 8421
rect 14461 8381 14473 8415
rect 14507 8381 14519 8415
rect 14642 8412 14648 8424
rect 14603 8384 14648 8412
rect 14461 8375 14519 8381
rect 12986 8344 12992 8356
rect 12406 8316 12992 8344
rect 12986 8304 12992 8316
rect 13044 8304 13050 8356
rect 14476 8344 14504 8375
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 17681 8415 17739 8421
rect 14752 8384 17632 8412
rect 14752 8344 14780 8384
rect 17034 8344 17040 8356
rect 14476 8316 14780 8344
rect 16995 8316 17040 8344
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 7834 8276 7840 8288
rect 7795 8248 7840 8276
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 9398 8236 9404 8288
rect 9456 8276 9462 8288
rect 9585 8279 9643 8285
rect 9585 8276 9597 8279
rect 9456 8248 9597 8276
rect 9456 8236 9462 8248
rect 9585 8245 9597 8248
rect 9631 8245 9643 8279
rect 17604 8276 17632 8384
rect 17681 8381 17693 8415
rect 17727 8381 17739 8415
rect 18506 8412 18512 8424
rect 18467 8384 18512 8412
rect 17681 8375 17739 8381
rect 17696 8344 17724 8375
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 19628 8412 19656 8520
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20671 8452 21404 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 18739 8384 19656 8412
rect 20088 8412 20116 8443
rect 20088 8384 21036 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 19518 8344 19524 8356
rect 17696 8316 19524 8344
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 21008 8353 21036 8384
rect 21376 8356 21404 8452
rect 20993 8347 21051 8353
rect 20993 8313 21005 8347
rect 21039 8344 21051 8347
rect 21174 8344 21180 8356
rect 21039 8316 21180 8344
rect 21039 8313 21051 8316
rect 20993 8307 21051 8313
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 21358 8344 21364 8356
rect 21319 8316 21364 8344
rect 21358 8304 21364 8316
rect 21416 8304 21422 8356
rect 17954 8276 17960 8288
rect 17604 8248 17960 8276
rect 9585 8239 9643 8245
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 9122 8072 9128 8084
rect 8343 8044 9128 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 10686 8072 10692 8084
rect 10647 8044 10692 8072
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 14424 8044 17049 8072
rect 14424 8032 14430 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 18932 8044 19349 8072
rect 18932 8032 18938 8044
rect 19337 8041 19349 8044
rect 19383 8041 19395 8075
rect 19337 8035 19395 8041
rect 10410 8004 10416 8016
rect 7668 7976 10416 8004
rect 7668 7945 7696 7976
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 16761 8007 16819 8013
rect 16761 7973 16773 8007
rect 16807 8004 16819 8007
rect 16942 8004 16948 8016
rect 16807 7976 16948 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 16942 7964 16948 7976
rect 17000 8004 17006 8016
rect 18506 8004 18512 8016
rect 17000 7976 18512 8004
rect 17000 7964 17006 7976
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7905 7711 7939
rect 7834 7936 7840 7948
rect 7795 7908 7840 7936
rect 7653 7899 7711 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 17512 7945 17540 7976
rect 18506 7964 18512 7976
rect 18564 7964 18570 8016
rect 12161 7939 12219 7945
rect 12161 7936 12173 7939
rect 11940 7908 12173 7936
rect 11940 7896 11946 7908
rect 12161 7905 12173 7908
rect 12207 7905 12219 7939
rect 12161 7899 12219 7905
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17678 7936 17684 7948
rect 17639 7908 17684 7936
rect 17497 7899 17555 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 18046 7936 18052 7948
rect 18007 7908 18052 7936
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 9398 7868 9404 7880
rect 9359 7840 9404 7868
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 13814 7868 13820 7880
rect 9723 7840 13820 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 20947 7840 21312 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 17405 7803 17463 7809
rect 17405 7769 17417 7803
rect 17451 7800 17463 7803
rect 17954 7800 17960 7812
rect 17451 7772 17960 7800
rect 17451 7769 17463 7772
rect 17405 7763 17463 7769
rect 17954 7760 17960 7772
rect 18012 7760 18018 7812
rect 21284 7744 21312 7840
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8202 7732 8208 7744
rect 7975 7704 8208 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 14976 7704 20729 7732
rect 14976 7692 14982 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 21266 7732 21272 7744
rect 21227 7704 21272 7732
rect 20717 7695 20775 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 7742 7528 7748 7540
rect 7703 7500 7748 7528
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8202 7528 8208 7540
rect 8163 7500 8208 7528
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 13630 7528 13636 7540
rect 9640 7500 13636 7528
rect 9640 7488 9646 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14645 7531 14703 7537
rect 14645 7497 14657 7531
rect 14691 7528 14703 7531
rect 18414 7528 18420 7540
rect 14691 7500 18420 7528
rect 14691 7497 14703 7500
rect 14645 7491 14703 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20346 7528 20352 7540
rect 20211 7500 20352 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 7760 7392 7788 7488
rect 7837 7463 7895 7469
rect 7837 7429 7849 7463
rect 7883 7460 7895 7463
rect 8294 7460 8300 7472
rect 7883 7432 8300 7460
rect 7883 7429 7895 7432
rect 7837 7423 7895 7429
rect 8294 7420 8300 7432
rect 8352 7460 8358 7472
rect 8849 7463 8907 7469
rect 8849 7460 8861 7463
rect 8352 7432 8861 7460
rect 8352 7420 8358 7432
rect 8849 7429 8861 7432
rect 8895 7460 8907 7463
rect 9398 7460 9404 7472
rect 8895 7432 9404 7460
rect 8895 7429 8907 7432
rect 8849 7423 8907 7429
rect 9398 7420 9404 7432
rect 9456 7420 9462 7472
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 19337 7463 19395 7469
rect 9548 7432 19104 7460
rect 9548 7420 9554 7432
rect 8478 7392 8484 7404
rect 7760 7364 8484 7392
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 10502 7392 10508 7404
rect 10463 7364 10508 7392
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 19076 7401 19104 7432
rect 19337 7429 19349 7463
rect 19383 7460 19395 7463
rect 20530 7460 20536 7472
rect 19383 7432 20536 7460
rect 19383 7429 19395 7432
rect 19337 7423 19395 7429
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 11348 7364 14473 7392
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 7340 7296 7573 7324
rect 7340 7284 7346 7296
rect 7561 7293 7573 7296
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 10321 7327 10379 7333
rect 10321 7293 10333 7327
rect 10367 7324 10379 7327
rect 11348 7324 11376 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 21082 7392 21088 7404
rect 21043 7364 21088 7392
rect 19981 7355 20039 7361
rect 11514 7324 11520 7336
rect 10367 7296 11376 7324
rect 11475 7296 11520 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 17954 7324 17960 7336
rect 17915 7296 17960 7324
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 19996 7324 20024 7355
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 18104 7296 20024 7324
rect 18104 7284 18110 7296
rect 17126 7216 17132 7268
rect 17184 7256 17190 7268
rect 20901 7259 20959 7265
rect 20901 7256 20913 7259
rect 17184 7228 20913 7256
rect 17184 7216 17190 7228
rect 20901 7225 20913 7228
rect 20947 7225 20959 7259
rect 20901 7219 20959 7225
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 15470 6984 15476 6996
rect 10744 6956 15476 6984
rect 10744 6944 10750 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 9582 6916 9588 6928
rect 8036 6888 9588 6916
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 8036 6857 8064 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 11146 6916 11152 6928
rect 11072 6888 11152 6916
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 1636 6820 7481 6848
rect 1636 6808 1642 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6848 9183 6851
rect 11072 6848 11100 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 9171 6820 11100 6848
rect 11164 6820 11437 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 7484 6780 7512 6811
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7484 6752 8125 6780
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9456 6752 10057 6780
rect 9456 6740 9462 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 11164 6780 11192 6820
rect 11425 6817 11437 6820
rect 11471 6848 11483 6851
rect 11790 6848 11796 6860
rect 11471 6820 11796 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6848 15255 6851
rect 17402 6848 17408 6860
rect 15243 6820 17408 6848
rect 15243 6817 15255 6820
rect 15197 6811 15255 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 10652 6752 11192 6780
rect 11241 6783 11299 6789
rect 10652 6740 10658 6752
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11514 6780 11520 6792
rect 11287 6752 11520 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 13228 6752 14289 6780
rect 13228 6740 13234 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 14599 6752 19257 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6780 20131 6783
rect 21085 6783 21143 6789
rect 20119 6752 20484 6780
rect 20119 6749 20131 6752
rect 20073 6743 20131 6749
rect 14642 6712 14648 6724
rect 9692 6684 14648 6712
rect 8202 6644 8208 6656
rect 8163 6616 8208 6644
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 8619 6616 9229 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 9217 6613 9229 6616
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9692 6653 9720 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 20456 6656 20484 6752
rect 21085 6749 21097 6783
rect 21131 6780 21143 6783
rect 21266 6780 21272 6792
rect 21131 6752 21272 6780
rect 21131 6749 21143 6752
rect 21085 6743 21143 6749
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 9677 6647 9735 6653
rect 9364 6616 9409 6644
rect 9364 6604 9370 6616
rect 9677 6613 9689 6647
rect 9723 6613 9735 6647
rect 9677 6607 9735 6613
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10836 6616 10885 6644
rect 10836 6604 10842 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 11885 6647 11943 6653
rect 11885 6644 11897 6647
rect 11379 6616 11897 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11885 6613 11897 6616
rect 11931 6644 11943 6647
rect 12526 6644 12532 6656
rect 11931 6616 12532 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 15286 6644 15292 6656
rect 15247 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15378 6604 15384 6656
rect 15436 6644 15442 6656
rect 15749 6647 15807 6653
rect 15436 6616 15481 6644
rect 15436 6604 15442 6616
rect 15749 6613 15761 6647
rect 15795 6644 15807 6647
rect 15930 6644 15936 6656
rect 15795 6616 15936 6644
rect 15795 6613 15807 6616
rect 15749 6607 15807 6613
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 19610 6644 19616 6656
rect 19475 6616 19616 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 19610 6604 19616 6616
rect 19668 6604 19674 6656
rect 19886 6644 19892 6656
rect 19847 6616 19892 6644
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 20438 6644 20444 6656
rect 20399 6616 20444 6644
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 20901 6647 20959 6653
rect 20901 6644 20913 6647
rect 20864 6616 20913 6644
rect 20864 6604 20870 6616
rect 20901 6613 20913 6616
rect 20947 6613 20959 6647
rect 20901 6607 20959 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 9217 6443 9275 6449
rect 9217 6409 9229 6443
rect 9263 6440 9275 6443
rect 9306 6440 9312 6452
rect 9263 6412 9312 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9456 6412 9597 6440
rect 9456 6400 9462 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10502 6440 10508 6452
rect 10459 6412 10508 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 9600 6372 9628 6403
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10778 6440 10784 6452
rect 10739 6412 10784 6440
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 13872 6412 14289 6440
rect 13872 6400 13878 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 14277 6403 14335 6409
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 15378 6440 15384 6452
rect 14783 6412 15384 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 17368 6412 20821 6440
rect 17368 6400 17374 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 20809 6403 20867 6409
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 21140 6412 21281 6440
rect 21140 6400 21146 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21269 6403 21327 6409
rect 16390 6372 16396 6384
rect 9600 6344 16396 6372
rect 16390 6332 16396 6344
rect 16448 6332 16454 6384
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 9490 6304 9496 6316
rect 8536 6276 9496 6304
rect 8536 6264 8542 6276
rect 9490 6264 9496 6276
rect 9548 6304 9554 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9548 6276 9689 6304
rect 9548 6264 9554 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11146 6304 11152 6316
rect 10919 6276 11152 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11756 6276 11897 6304
rect 11756 6264 11762 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 14369 6307 14427 6313
rect 12032 6276 13952 6304
rect 12032 6264 12038 6276
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6205 9827 6239
rect 11054 6236 11060 6248
rect 11015 6208 11060 6236
rect 9769 6199 9827 6205
rect 9582 6128 9588 6180
rect 9640 6168 9646 6180
rect 9784 6168 9812 6199
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6205 11667 6239
rect 11609 6199 11667 6205
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12526 6236 12532 6248
rect 11839 6208 12532 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 9640 6140 9812 6168
rect 11624 6168 11652 6199
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12434 6168 12440 6180
rect 11624 6140 12440 6168
rect 9640 6128 9646 6140
rect 12434 6128 12440 6140
rect 12492 6168 12498 6180
rect 13630 6168 13636 6180
rect 12492 6140 13636 6168
rect 12492 6128 12498 6140
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 13924 6168 13952 6276
rect 14108 6276 14320 6304
rect 14108 6245 14136 6276
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6205 14151 6239
rect 14292 6236 14320 6276
rect 14369 6273 14381 6307
rect 14415 6304 14427 6307
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14415 6276 15025 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 19058 6264 19064 6316
rect 19116 6304 19122 6316
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 19116 6276 20453 6304
rect 19116 6264 19122 6276
rect 20441 6273 20453 6276
rect 20487 6304 20499 6307
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 20487 6276 21005 6304
rect 20487 6273 20499 6276
rect 20441 6267 20499 6273
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 16022 6236 16028 6248
rect 14292 6208 16028 6236
rect 14093 6199 14151 6205
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 15378 6168 15384 6180
rect 13924 6140 15384 6168
rect 15378 6128 15384 6140
rect 15436 6128 15442 6180
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8260 6072 8769 6100
rect 8260 6060 8266 6072
rect 8757 6069 8769 6072
rect 8803 6100 8815 6103
rect 11974 6100 11980 6112
rect 8803 6072 11980 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12526 6100 12532 6112
rect 12487 6072 12532 6100
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 9548 5868 10241 5896
rect 9548 5856 9554 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 10229 5859 10287 5865
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 13096 5828 13124 5859
rect 13096 5800 14136 5828
rect 11698 5760 11704 5772
rect 11659 5732 11704 5760
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 13078 5760 13084 5772
rect 12575 5732 13084 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 14108 5701 14136 5800
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5760 14427 5763
rect 18046 5760 18052 5772
rect 14415 5732 18052 5760
rect 14415 5729 14427 5732
rect 14369 5723 14427 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12308 5664 12725 5692
rect 12308 5652 12314 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 15010 5624 15016 5636
rect 4120 5596 15016 5624
rect 4120 5584 4126 5596
rect 15010 5584 15016 5596
rect 15068 5584 15074 5636
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 12434 5556 12440 5568
rect 9548 5528 12440 5556
rect 9548 5516 9554 5528
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 21266 5556 21272 5568
rect 21227 5528 21272 5556
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 1486 5312 1492 5364
rect 1544 5352 1550 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 1544 5324 8309 5352
rect 1544 5312 1550 5324
rect 8297 5321 8309 5324
rect 8343 5352 8355 5355
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8343 5324 8953 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 8941 5315 8999 5321
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 13081 5355 13139 5361
rect 13081 5352 13093 5355
rect 12676 5324 13093 5352
rect 12676 5312 12682 5324
rect 13081 5321 13093 5324
rect 13127 5321 13139 5355
rect 15286 5352 15292 5364
rect 15247 5324 15292 5352
rect 13081 5315 13139 5321
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 18138 5352 18144 5364
rect 15620 5324 18144 5352
rect 15620 5312 15626 5324
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 13449 5287 13507 5293
rect 13449 5284 13461 5287
rect 11072 5256 13461 5284
rect 11072 5228 11100 5256
rect 13449 5253 13461 5256
rect 13495 5284 13507 5287
rect 14093 5287 14151 5293
rect 14093 5284 14105 5287
rect 13495 5256 14105 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 14093 5253 14105 5256
rect 14139 5253 14151 5287
rect 14093 5247 14151 5253
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5216 9091 5219
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9079 5188 9689 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9677 5185 9689 5188
rect 9723 5216 9735 5219
rect 11054 5216 11060 5228
rect 9723 5188 11060 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 12710 5216 12716 5228
rect 12671 5188 12716 5216
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9490 5148 9496 5160
rect 8895 5120 9496 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 12728 5148 12756 5176
rect 13541 5151 13599 5157
rect 13541 5148 13553 5151
rect 12728 5120 13553 5148
rect 13541 5117 13553 5120
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 15746 5148 15752 5160
rect 13688 5120 13733 5148
rect 15707 5120 15752 5148
rect 13688 5108 13694 5120
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 16022 5148 16028 5160
rect 15979 5120 16028 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 18690 5080 18696 5092
rect 12268 5052 18696 5080
rect 12268 5024 12296 5052
rect 18690 5040 18696 5052
rect 18748 5040 18754 5092
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 9272 4984 9413 5012
rect 9272 4972 9278 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 9401 4975 9459 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 12250 5012 12256 5024
rect 12211 4984 12256 5012
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 13170 4808 13176 4820
rect 9723 4780 12756 4808
rect 13131 4780 13176 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4641 9091 4675
rect 9214 4672 9220 4684
rect 9175 4644 9220 4672
rect 9033 4635 9091 4641
rect 9048 4604 9076 4635
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 9548 4644 10609 4672
rect 9548 4632 9554 4644
rect 10597 4641 10609 4644
rect 10643 4672 10655 4675
rect 10686 4672 10692 4684
rect 10643 4644 10692 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 11517 4675 11575 4681
rect 11517 4641 11529 4675
rect 11563 4672 11575 4675
rect 12250 4672 12256 4684
rect 11563 4644 12256 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9048 4576 9965 4604
rect 9953 4573 9965 4576
rect 9999 4604 10011 4607
rect 11532 4604 11560 4635
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12728 4681 12756 4780
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 12713 4675 12771 4681
rect 12713 4641 12725 4675
rect 12759 4641 12771 4675
rect 12713 4635 12771 4641
rect 9999 4576 11560 4604
rect 12636 4604 12664 4635
rect 14734 4604 14740 4616
rect 12636 4576 14740 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 10689 4539 10747 4545
rect 10689 4536 10701 4539
rect 8444 4508 10701 4536
rect 8444 4496 8450 4508
rect 10689 4505 10701 4508
rect 10735 4536 10747 4539
rect 11514 4536 11520 4548
rect 10735 4508 11520 4536
rect 10735 4505 10747 4508
rect 10689 4499 10747 4505
rect 11514 4496 11520 4508
rect 11572 4536 11578 4548
rect 11882 4536 11888 4548
rect 11572 4508 11888 4536
rect 11572 4496 11578 4508
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 12805 4539 12863 4545
rect 12805 4536 12817 4539
rect 12406 4508 12817 4536
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 9364 4440 9409 4468
rect 9364 4428 9370 4440
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 11149 4471 11207 4477
rect 10836 4440 10881 4468
rect 10836 4428 10842 4440
rect 11149 4437 11161 4471
rect 11195 4468 11207 4471
rect 11701 4471 11759 4477
rect 11701 4468 11713 4471
rect 11195 4440 11713 4468
rect 11195 4437 11207 4440
rect 11149 4431 11207 4437
rect 11701 4437 11713 4440
rect 11747 4437 11759 4471
rect 11701 4431 11759 4437
rect 11793 4471 11851 4477
rect 11793 4437 11805 4471
rect 11839 4468 11851 4471
rect 12066 4468 12072 4480
rect 11839 4440 12072 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12161 4471 12219 4477
rect 12161 4437 12173 4471
rect 12207 4468 12219 4471
rect 12406 4468 12434 4508
rect 12805 4505 12817 4508
rect 12851 4505 12863 4539
rect 12805 4499 12863 4505
rect 12207 4440 12434 4468
rect 12207 4437 12219 4440
rect 12161 4431 12219 4437
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 9217 4267 9275 4273
rect 9217 4233 9229 4267
rect 9263 4264 9275 4267
rect 9306 4264 9312 4276
rect 9263 4236 9312 4264
rect 9263 4233 9275 4236
rect 9217 4227 9275 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9585 4267 9643 4273
rect 9585 4233 9597 4267
rect 9631 4264 9643 4267
rect 10042 4264 10048 4276
rect 9631 4236 10048 4264
rect 9631 4233 9643 4236
rect 9585 4227 9643 4233
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 10836 4236 11529 4264
rect 10836 4224 10842 4236
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 12066 4264 12072 4276
rect 12027 4236 12072 4264
rect 11517 4227 11575 4233
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 11054 4196 11060 4208
rect 9548 4168 9812 4196
rect 9548 4156 9554 4168
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 1452 4032 2774 4060
rect 1452 4020 1458 4032
rect 2746 3992 2774 4032
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9490 4060 9496 4072
rect 8720 4032 9496 4060
rect 8720 4020 8726 4032
rect 9490 4020 9496 4032
rect 9548 4060 9554 4072
rect 9784 4069 9812 4168
rect 10796 4168 11060 4196
rect 10594 4128 10600 4140
rect 10520 4100 10600 4128
rect 10520 4069 10548 4100
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10796 4137 10824 4168
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 11532 4196 11560 4227
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 12526 4264 12532 4276
rect 12406 4236 12532 4264
rect 12406 4196 12434 4236
rect 12526 4224 12532 4236
rect 12584 4264 12590 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 12584 4236 13461 4264
rect 12584 4224 12590 4236
rect 13449 4233 13461 4236
rect 13495 4264 13507 4267
rect 14553 4267 14611 4273
rect 14553 4264 14565 4267
rect 13495 4236 14565 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 14553 4233 14565 4236
rect 14599 4264 14611 4267
rect 17954 4264 17960 4276
rect 14599 4236 17960 4264
rect 14599 4233 14611 4236
rect 14553 4227 14611 4233
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 11532 4168 12434 4196
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 13188 4100 13400 4128
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9548 4032 9689 4060
rect 9548 4020 9554 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 10594 3992 10600 4004
rect 2746 3964 10600 3992
rect 10594 3952 10600 3964
rect 10652 3992 10658 4004
rect 10704 3992 10732 4023
rect 11146 3992 11152 4004
rect 10652 3964 10732 3992
rect 11107 3964 11152 3992
rect 10652 3952 10658 3964
rect 11146 3952 11152 3964
rect 11204 3952 11210 4004
rect 11882 3952 11888 4004
rect 11940 3992 11946 4004
rect 13188 3992 13216 4100
rect 13372 4069 13400 4100
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 18046 4128 18052 4140
rect 16448 4100 18052 4128
rect 16448 4088 16454 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 13403 4032 14197 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 14185 4029 14197 4032
rect 14231 4060 14243 4063
rect 17954 4060 17960 4072
rect 14231 4032 17960 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 11940 3964 13216 3992
rect 11940 3952 11946 3964
rect 13280 3924 13308 4023
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 13814 3992 13820 4004
rect 13775 3964 13820 3992
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 15289 3995 15347 4001
rect 15289 3992 15301 3995
rect 14608 3964 15301 3992
rect 14608 3952 14614 3964
rect 15289 3961 15301 3964
rect 15335 3992 15347 3995
rect 18966 3992 18972 4004
rect 15335 3964 18972 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 18966 3952 18972 3964
rect 19024 3952 19030 4004
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 13280 3896 14933 3924
rect 14921 3893 14933 3896
rect 14967 3924 14979 3927
rect 15470 3924 15476 3936
rect 14967 3896 15476 3924
rect 14967 3893 14979 3896
rect 14921 3887 14979 3893
rect 15470 3884 15476 3896
rect 15528 3924 15534 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15528 3896 15669 3924
rect 15528 3884 15534 3896
rect 15657 3893 15669 3896
rect 15703 3924 15715 3927
rect 17586 3924 17592 3936
rect 15703 3896 17592 3924
rect 15703 3893 15715 3896
rect 15657 3887 15715 3893
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 9548 3692 9873 3720
rect 9548 3680 9554 3692
rect 9861 3689 9873 3692
rect 9907 3689 9919 3723
rect 9861 3683 9919 3689
rect 9876 3380 9904 3683
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10100 3692 10241 3720
rect 10100 3680 10106 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10594 3720 10600 3732
rect 10555 3692 10600 3720
rect 10229 3683 10287 3689
rect 10244 3448 10272 3683
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 11112 3692 11253 3720
rect 11112 3680 11118 3692
rect 11241 3689 11253 3692
rect 11287 3720 11299 3723
rect 15013 3723 15071 3729
rect 11287 3692 12434 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 12406 3516 12434 3692
rect 15013 3689 15025 3723
rect 15059 3720 15071 3723
rect 15654 3720 15660 3732
rect 15059 3692 15660 3720
rect 15059 3689 15071 3692
rect 15013 3683 15071 3689
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 16025 3723 16083 3729
rect 16025 3720 16037 3723
rect 15804 3692 16037 3720
rect 15804 3680 15810 3692
rect 16025 3689 16037 3692
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 17129 3723 17187 3729
rect 17129 3689 17141 3723
rect 17175 3720 17187 3723
rect 17586 3720 17592 3732
rect 17175 3692 17592 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 14384 3624 15516 3652
rect 14384 3593 14412 3624
rect 15488 3596 15516 3624
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3553 14427 3587
rect 14550 3584 14556 3596
rect 14511 3556 14556 3584
rect 14369 3547 14427 3553
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3584 16543 3587
rect 17770 3584 17776 3596
rect 16531 3556 17776 3584
rect 16531 3553 16543 3556
rect 16485 3547 16543 3553
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 16761 3519 16819 3525
rect 12406 3488 15700 3516
rect 10244 3420 14688 3448
rect 14660 3392 14688 3420
rect 15672 3392 15700 3488
rect 16761 3485 16773 3519
rect 16807 3516 16819 3519
rect 17034 3516 17040 3528
rect 16807 3488 17040 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 14550 3380 14556 3392
rect 9876 3352 14556 3380
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 15562 3380 15568 3392
rect 14700 3352 14745 3380
rect 15523 3352 15568 3380
rect 14700 3340 14706 3352
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 15712 3352 15757 3380
rect 15712 3340 15718 3352
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 15197 3179 15255 3185
rect 15197 3176 15209 3179
rect 12216 3148 15209 3176
rect 12216 3136 12222 3148
rect 15197 3145 15209 3148
rect 15243 3176 15255 3179
rect 15562 3176 15568 3188
rect 15243 3148 15568 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 14700 3012 15577 3040
rect 14700 3000 14706 3012
rect 15565 3009 15577 3012
rect 15611 3040 15623 3043
rect 17954 3040 17960 3052
rect 15611 3012 17960 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 16209 2839 16267 2845
rect 16209 2836 16221 2839
rect 15712 2808 16221 2836
rect 15712 2796 15718 2808
rect 16209 2805 16221 2808
rect 16255 2836 16267 2839
rect 19058 2836 19064 2848
rect 16255 2808 19064 2836
rect 16255 2805 16267 2808
rect 16209 2799 16267 2805
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 19150 2632 19156 2644
rect 15436 2604 19156 2632
rect 15436 2592 15442 2604
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 19242 2564 19248 2576
rect 12492 2536 19248 2564
rect 12492 2524 12498 2536
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 13084 20544 13136 20596
rect 20628 20544 20680 20596
rect 21548 20544 21600 20596
rect 7288 20476 7340 20528
rect 10600 20408 10652 20460
rect 9312 20340 9364 20392
rect 17316 20340 17368 20392
rect 5724 20272 5776 20324
rect 19616 20272 19668 20324
rect 18144 20204 18196 20256
rect 18788 20247 18840 20256
rect 18788 20213 18797 20247
rect 18797 20213 18831 20247
rect 18831 20213 18840 20247
rect 18788 20204 18840 20213
rect 18880 20204 18932 20256
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 5724 20043 5776 20052
rect 5724 20009 5733 20043
rect 5733 20009 5767 20043
rect 5767 20009 5776 20043
rect 5724 20000 5776 20009
rect 11980 20000 12032 20052
rect 17868 20000 17920 20052
rect 18604 20000 18656 20052
rect 20260 20000 20312 20052
rect 4160 19839 4212 19848
rect 4160 19805 4169 19839
rect 4169 19805 4203 19839
rect 4203 19805 4212 19839
rect 4160 19796 4212 19805
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 9128 19864 9180 19916
rect 9312 19864 9364 19916
rect 12256 19864 12308 19916
rect 17960 19932 18012 19984
rect 19708 19932 19760 19984
rect 20812 19932 20864 19984
rect 19248 19864 19300 19916
rect 21272 19864 21324 19916
rect 4344 19703 4396 19712
rect 4344 19669 4353 19703
rect 4353 19669 4387 19703
rect 4387 19669 4396 19703
rect 4344 19660 4396 19669
rect 11244 19796 11296 19848
rect 11704 19796 11756 19848
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 17132 19796 17184 19848
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 17776 19796 17828 19848
rect 18236 19796 18288 19848
rect 18788 19796 18840 19848
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 20260 19796 20312 19848
rect 20628 19796 20680 19848
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 18420 19728 18472 19780
rect 17684 19660 17736 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 13728 19456 13780 19508
rect 21364 19456 21416 19508
rect 1400 19388 1452 19440
rect 2596 19388 2648 19440
rect 4252 19388 4304 19440
rect 4804 19388 4856 19440
rect 7288 19431 7340 19440
rect 7288 19397 7297 19431
rect 7297 19397 7331 19431
rect 7331 19397 7340 19431
rect 7288 19388 7340 19397
rect 4528 19320 4580 19372
rect 7564 19363 7616 19372
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 11704 19388 11756 19440
rect 12900 19388 12952 19440
rect 15384 19388 15436 19440
rect 16396 19388 16448 19440
rect 10784 19320 10836 19372
rect 11520 19320 11572 19372
rect 14372 19320 14424 19372
rect 17868 19388 17920 19440
rect 20996 19388 21048 19440
rect 22468 19388 22520 19440
rect 3976 19252 4028 19304
rect 6644 19252 6696 19304
rect 9772 19252 9824 19304
rect 10876 19252 10928 19304
rect 13268 19252 13320 19304
rect 16948 19252 17000 19304
rect 18512 19320 18564 19372
rect 21180 19320 21232 19372
rect 940 19184 992 19236
rect 5816 19184 5868 19236
rect 4344 19116 4396 19168
rect 11520 19159 11572 19168
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 13268 19159 13320 19168
rect 13268 19125 13277 19159
rect 13277 19125 13311 19159
rect 13311 19125 13320 19159
rect 13268 19116 13320 19125
rect 13728 19116 13780 19168
rect 19524 19184 19576 19236
rect 20444 19184 20496 19236
rect 18604 19116 18656 19168
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 19064 19159 19116 19168
rect 18696 19116 18748 19125
rect 19064 19125 19073 19159
rect 19073 19125 19107 19159
rect 19107 19125 19116 19159
rect 19064 19116 19116 19125
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 3148 18912 3200 18964
rect 7380 18912 7432 18964
rect 16304 18955 16356 18964
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 5172 18751 5224 18760
rect 4160 18640 4212 18692
rect 4896 18683 4948 18692
rect 4896 18649 4905 18683
rect 4905 18649 4939 18683
rect 4939 18649 4948 18683
rect 4896 18640 4948 18649
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 7748 18640 7800 18692
rect 16304 18921 16313 18955
rect 16313 18921 16347 18955
rect 16347 18921 16356 18955
rect 16304 18912 16356 18921
rect 9128 18819 9180 18828
rect 9128 18785 9137 18819
rect 9137 18785 9171 18819
rect 9171 18785 9180 18819
rect 9128 18776 9180 18785
rect 8668 18708 8720 18760
rect 9036 18708 9088 18760
rect 12440 18708 12492 18760
rect 13728 18708 13780 18760
rect 17868 18708 17920 18760
rect 19064 18708 19116 18760
rect 21272 18708 21324 18760
rect 11060 18640 11112 18692
rect 11152 18640 11204 18692
rect 11980 18640 12032 18692
rect 13176 18640 13228 18692
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 10692 18615 10744 18624
rect 10692 18581 10701 18615
rect 10701 18581 10735 18615
rect 10735 18581 10744 18615
rect 10692 18572 10744 18581
rect 11704 18572 11756 18624
rect 13636 18572 13688 18624
rect 15476 18640 15528 18692
rect 17132 18640 17184 18692
rect 17500 18640 17552 18692
rect 19524 18640 19576 18692
rect 16304 18572 16356 18624
rect 16948 18572 17000 18624
rect 17316 18615 17368 18624
rect 17316 18581 17325 18615
rect 17325 18581 17359 18615
rect 17359 18581 17368 18615
rect 17316 18572 17368 18581
rect 21180 18572 21232 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 388 18368 440 18420
rect 6460 18368 6512 18420
rect 8668 18411 8720 18420
rect 8668 18377 8677 18411
rect 8677 18377 8711 18411
rect 8711 18377 8720 18411
rect 8668 18368 8720 18377
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 12440 18368 12492 18420
rect 12532 18368 12584 18420
rect 12716 18368 12768 18420
rect 13728 18368 13780 18420
rect 16948 18368 17000 18420
rect 17408 18368 17460 18420
rect 18972 18368 19024 18420
rect 4528 18343 4580 18352
rect 4528 18309 4537 18343
rect 4537 18309 4571 18343
rect 4571 18309 4580 18343
rect 4528 18300 4580 18309
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 10692 18300 10744 18352
rect 11060 18300 11112 18352
rect 15200 18300 15252 18352
rect 7748 18232 7800 18284
rect 8668 18232 8720 18284
rect 10968 18232 11020 18284
rect 13636 18232 13688 18284
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 9312 18164 9364 18216
rect 20904 18300 20956 18352
rect 21180 18300 21232 18352
rect 18144 18232 18196 18284
rect 18696 18232 18748 18284
rect 21456 18232 21508 18284
rect 4896 18096 4948 18148
rect 11704 18096 11756 18148
rect 6552 18028 6604 18080
rect 6920 18028 6972 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 9496 18028 9548 18080
rect 12348 18071 12400 18080
rect 12348 18037 12357 18071
rect 12357 18037 12391 18071
rect 12391 18037 12400 18071
rect 12348 18028 12400 18037
rect 17868 18164 17920 18216
rect 14280 18096 14332 18148
rect 17500 18096 17552 18148
rect 13820 18028 13872 18080
rect 15292 18028 15344 18080
rect 19524 18028 19576 18080
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 4712 17824 4764 17876
rect 5908 17824 5960 17876
rect 3884 17731 3936 17740
rect 3884 17697 3893 17731
rect 3893 17697 3927 17731
rect 3927 17697 3936 17731
rect 3884 17688 3936 17697
rect 9588 17756 9640 17808
rect 10232 17824 10284 17876
rect 13176 17867 13228 17876
rect 5632 17731 5684 17740
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 9220 17731 9272 17740
rect 6000 17620 6052 17672
rect 9220 17697 9229 17731
rect 9229 17697 9263 17731
rect 9263 17697 9272 17731
rect 9220 17688 9272 17697
rect 10324 17688 10376 17740
rect 4344 17484 4396 17536
rect 7196 17552 7248 17604
rect 8484 17552 8536 17604
rect 9588 17484 9640 17536
rect 9680 17484 9732 17536
rect 10508 17484 10560 17536
rect 12440 17620 12492 17672
rect 10692 17552 10744 17604
rect 13176 17833 13185 17867
rect 13185 17833 13219 17867
rect 13219 17833 13228 17867
rect 13176 17824 13228 17833
rect 13728 17824 13780 17876
rect 17868 17824 17920 17876
rect 13084 17620 13136 17672
rect 17316 17620 17368 17672
rect 20904 17663 20956 17672
rect 20904 17629 20922 17663
rect 20922 17629 20956 17663
rect 20904 17620 20956 17629
rect 21272 17620 21324 17672
rect 18144 17552 18196 17604
rect 19708 17484 19760 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 4344 17323 4396 17332
rect 4344 17289 4353 17323
rect 4353 17289 4387 17323
rect 4387 17289 4396 17323
rect 4344 17280 4396 17289
rect 4804 17280 4856 17332
rect 5632 17280 5684 17332
rect 7840 17212 7892 17264
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 10416 17280 10468 17332
rect 12440 17212 12492 17264
rect 15752 17255 15804 17264
rect 11612 17144 11664 17196
rect 11796 17187 11848 17196
rect 11796 17153 11830 17187
rect 11830 17153 11848 17187
rect 11796 17144 11848 17153
rect 12348 17144 12400 17196
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 9680 17008 9732 17060
rect 11152 17008 11204 17060
rect 13084 17008 13136 17060
rect 12992 16940 13044 16992
rect 15752 17221 15761 17255
rect 15761 17221 15795 17255
rect 15795 17221 15804 17255
rect 15752 17212 15804 17221
rect 14372 17187 14424 17196
rect 14372 17153 14406 17187
rect 14406 17153 14424 17187
rect 14372 17144 14424 17153
rect 17868 17280 17920 17332
rect 19708 17144 19760 17196
rect 15200 16940 15252 16992
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 6828 16736 6880 16788
rect 6920 16736 6972 16788
rect 4528 16643 4580 16652
rect 4528 16609 4537 16643
rect 4537 16609 4571 16643
rect 4571 16609 4580 16643
rect 4528 16600 4580 16609
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 9220 16736 9272 16788
rect 12348 16736 12400 16788
rect 9496 16600 9548 16652
rect 10968 16600 11020 16652
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 15476 16736 15528 16788
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 15200 16575 15252 16584
rect 6000 16464 6052 16516
rect 7288 16464 7340 16516
rect 2412 16396 2464 16448
rect 5540 16396 5592 16448
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7840 16439 7892 16448
rect 7196 16396 7248 16405
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 8668 16396 8720 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 15200 16541 15218 16575
rect 15218 16541 15252 16575
rect 15200 16532 15252 16541
rect 15752 16532 15804 16584
rect 17868 16600 17920 16652
rect 21272 16643 21324 16652
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 11704 16464 11756 16516
rect 15292 16464 15344 16516
rect 17592 16464 17644 16516
rect 12072 16396 12124 16448
rect 12532 16396 12584 16448
rect 12900 16396 12952 16448
rect 13452 16396 13504 16448
rect 13820 16396 13872 16448
rect 15200 16396 15252 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 5540 16192 5592 16244
rect 5724 16192 5776 16244
rect 6000 16124 6052 16176
rect 6736 16124 6788 16176
rect 10048 16192 10100 16244
rect 11980 16192 12032 16244
rect 12072 16192 12124 16244
rect 17592 16192 17644 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 8392 16056 8444 16108
rect 13176 16124 13228 16176
rect 12992 16099 13044 16108
rect 12992 16065 13010 16099
rect 13010 16065 13044 16099
rect 12992 16056 13044 16065
rect 20536 16056 20588 16108
rect 21272 16056 21324 16108
rect 8392 15852 8444 15904
rect 13452 15852 13504 15904
rect 14464 15852 14516 15904
rect 19064 15852 19116 15904
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 21272 15691 21324 15700
rect 21272 15657 21281 15691
rect 21281 15657 21315 15691
rect 21315 15657 21324 15691
rect 21272 15648 21324 15657
rect 14280 15512 14332 15564
rect 13452 15444 13504 15496
rect 17868 15444 17920 15496
rect 13176 15376 13228 15428
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 13452 15308 13504 15360
rect 18144 15376 18196 15428
rect 19524 15376 19576 15428
rect 17684 15308 17736 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 5172 15104 5224 15156
rect 6828 15104 6880 15156
rect 8116 15104 8168 15156
rect 7104 15036 7156 15088
rect 9956 15036 10008 15088
rect 16396 15036 16448 15088
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 7656 14968 7708 15020
rect 16212 15011 16264 15020
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 17868 15104 17920 15156
rect 20720 15036 20772 15088
rect 16212 14968 16264 14977
rect 21272 14968 21324 15020
rect 14372 14900 14424 14952
rect 15200 14832 15252 14884
rect 4528 14764 4580 14816
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 9680 14764 9732 14816
rect 12992 14764 13044 14816
rect 14280 14764 14332 14816
rect 19524 14764 19576 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 5632 14424 5684 14476
rect 9680 14492 9732 14544
rect 8208 14424 8260 14476
rect 11704 14560 11756 14612
rect 8116 14263 8168 14272
rect 8116 14229 8125 14263
rect 8125 14229 8159 14263
rect 8159 14229 8168 14263
rect 8116 14220 8168 14229
rect 9496 14220 9548 14272
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 12440 14356 12492 14408
rect 16212 14560 16264 14612
rect 19248 14560 19300 14612
rect 16396 14492 16448 14544
rect 21272 14560 21324 14612
rect 13084 14288 13136 14340
rect 10508 14220 10560 14272
rect 17316 14356 17368 14408
rect 19984 14356 20036 14408
rect 15200 14331 15252 14340
rect 15200 14297 15218 14331
rect 15218 14297 15252 14331
rect 15200 14288 15252 14297
rect 15476 14288 15528 14340
rect 13452 14220 13504 14272
rect 13728 14220 13780 14272
rect 20720 14263 20772 14272
rect 20720 14229 20729 14263
rect 20729 14229 20763 14263
rect 20763 14229 20772 14263
rect 20720 14220 20772 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 4252 14016 4304 14068
rect 8116 14016 8168 14068
rect 9312 14016 9364 14068
rect 9404 14016 9456 14068
rect 10692 14016 10744 14068
rect 15476 14016 15528 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 21272 14016 21324 14068
rect 13452 13948 13504 14000
rect 10048 13812 10100 13864
rect 11704 13812 11756 13864
rect 13452 13812 13504 13864
rect 16212 13812 16264 13864
rect 19340 13812 19392 13864
rect 20076 13812 20128 13864
rect 11888 13744 11940 13796
rect 9588 13676 9640 13728
rect 11612 13676 11664 13728
rect 16396 13744 16448 13796
rect 17592 13676 17644 13728
rect 19708 13676 19760 13728
rect 21180 13676 21232 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 4436 13472 4488 13524
rect 7288 13472 7340 13524
rect 7748 13472 7800 13524
rect 8024 13472 8076 13524
rect 9772 13472 9824 13524
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 13452 13515 13504 13524
rect 11612 13404 11664 13456
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 16212 13472 16264 13524
rect 18052 13472 18104 13524
rect 7288 13268 7340 13320
rect 10876 13268 10928 13320
rect 13452 13268 13504 13320
rect 17592 13268 17644 13320
rect 6736 13200 6788 13252
rect 8300 13200 8352 13252
rect 12440 13200 12492 13252
rect 13728 13200 13780 13252
rect 15568 13200 15620 13252
rect 18420 13268 18472 13320
rect 20812 13336 20864 13388
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 13360 13132 13412 13184
rect 13544 13132 13596 13184
rect 14832 13132 14884 13184
rect 16028 13132 16080 13184
rect 18052 13200 18104 13252
rect 19340 13132 19392 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 7564 12928 7616 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 13452 12971 13504 12980
rect 10508 12928 10560 12937
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 18420 12971 18472 12980
rect 18420 12937 18429 12971
rect 18429 12937 18463 12971
rect 18463 12937 18472 12971
rect 18420 12928 18472 12937
rect 11152 12860 11204 12912
rect 12532 12792 12584 12844
rect 20812 12860 20864 12912
rect 21272 12860 21324 12912
rect 15476 12724 15528 12776
rect 17684 12656 17736 12708
rect 9588 12588 9640 12640
rect 13820 12588 13872 12640
rect 15660 12588 15712 12640
rect 17960 12588 18012 12640
rect 18880 12588 18932 12640
rect 19248 12588 19300 12640
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 12348 12384 12400 12436
rect 16028 12384 16080 12436
rect 11244 12248 11296 12300
rect 10140 12180 10192 12232
rect 16948 12180 17000 12232
rect 17224 12180 17276 12232
rect 18420 12180 18472 12232
rect 19984 12180 20036 12232
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 12716 12112 12768 12164
rect 15200 12112 15252 12164
rect 15292 12112 15344 12164
rect 6736 12044 6788 12096
rect 6828 12044 6880 12096
rect 14280 12044 14332 12096
rect 16028 12044 16080 12096
rect 18420 12044 18472 12096
rect 18696 12044 18748 12096
rect 19800 12044 19852 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 6736 11883 6788 11892
rect 6736 11849 6745 11883
rect 6745 11849 6779 11883
rect 6779 11849 6788 11883
rect 6736 11840 6788 11849
rect 7012 11772 7064 11824
rect 12808 11840 12860 11892
rect 17040 11840 17092 11892
rect 14556 11772 14608 11824
rect 15200 11772 15252 11824
rect 19064 11840 19116 11892
rect 17868 11772 17920 11824
rect 13636 11704 13688 11756
rect 6828 11636 6880 11688
rect 11152 11568 11204 11620
rect 13360 11568 13412 11620
rect 7288 11500 7340 11552
rect 12808 11500 12860 11552
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 18420 11747 18472 11756
rect 18420 11713 18438 11747
rect 18438 11713 18472 11747
rect 18696 11772 18748 11824
rect 18420 11704 18472 11713
rect 19800 11704 19852 11756
rect 20904 11704 20956 11756
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 15016 11500 15068 11552
rect 17408 11500 17460 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 12900 11296 12952 11348
rect 13360 11296 13412 11348
rect 17684 11296 17736 11348
rect 20536 11296 20588 11348
rect 20904 11339 20956 11348
rect 20904 11305 20913 11339
rect 20913 11305 20947 11339
rect 20947 11305 20956 11339
rect 20904 11296 20956 11305
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 19064 11160 19116 11212
rect 11796 11024 11848 11076
rect 12348 11024 12400 11076
rect 13268 11092 13320 11144
rect 13452 11092 13504 11144
rect 17040 11135 17092 11144
rect 17040 11101 17058 11135
rect 17058 11101 17092 11135
rect 17316 11135 17368 11144
rect 17040 11092 17092 11101
rect 11060 10956 11112 11008
rect 12900 10956 12952 11008
rect 13544 10956 13596 11008
rect 13820 11024 13872 11076
rect 15016 11024 15068 11076
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 18696 11092 18748 11144
rect 19156 11024 19208 11076
rect 15200 10956 15252 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 8208 10752 8260 10804
rect 7380 10684 7432 10736
rect 7104 10616 7156 10668
rect 12900 10752 12952 10804
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 8116 10412 8168 10464
rect 8208 10412 8260 10464
rect 9404 10548 9456 10600
rect 11060 10548 11112 10600
rect 14740 10659 14792 10668
rect 14740 10625 14758 10659
rect 14758 10625 14792 10659
rect 14740 10616 14792 10625
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 17408 10752 17460 10804
rect 17316 10684 17368 10736
rect 15016 10616 15068 10625
rect 16856 10616 16908 10668
rect 19156 10752 19208 10804
rect 20904 10752 20956 10804
rect 21272 10616 21324 10668
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 15568 10412 15620 10464
rect 16488 10412 16540 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 12716 10208 12768 10260
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 15292 10208 15344 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 10600 10072 10652 10124
rect 17316 10072 17368 10124
rect 12256 10004 12308 10056
rect 12900 10004 12952 10056
rect 16488 10004 16540 10056
rect 11244 9868 11296 9920
rect 11704 9868 11756 9920
rect 15016 9868 15068 9920
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 9312 9664 9364 9716
rect 17224 9664 17276 9716
rect 6644 9596 6696 9648
rect 13820 9596 13872 9648
rect 7656 9528 7708 9580
rect 8668 9528 8720 9580
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 15108 9528 15160 9580
rect 20536 9571 20588 9580
rect 6552 9460 6604 9512
rect 5724 9392 5776 9444
rect 11244 9460 11296 9512
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 12348 9392 12400 9444
rect 14464 9392 14516 9444
rect 15660 9435 15712 9444
rect 15660 9401 15669 9435
rect 15669 9401 15703 9435
rect 15703 9401 15712 9435
rect 15660 9392 15712 9401
rect 19892 9435 19944 9444
rect 19892 9401 19901 9435
rect 19901 9401 19935 9435
rect 19935 9401 19944 9435
rect 19892 9392 19944 9401
rect 20628 9392 20680 9444
rect 12716 9324 12768 9376
rect 17132 9324 17184 9376
rect 21180 9367 21232 9376
rect 21180 9333 21189 9367
rect 21189 9333 21223 9367
rect 21223 9333 21232 9367
rect 21180 9324 21232 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 10692 9120 10744 9172
rect 12348 9120 12400 9172
rect 14188 9163 14240 9172
rect 14188 9129 14197 9163
rect 14197 9129 14231 9163
rect 14231 9129 14240 9163
rect 14188 9120 14240 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 17224 9163 17276 9172
rect 15292 9120 15344 9129
rect 17224 9129 17233 9163
rect 17233 9129 17267 9163
rect 17267 9129 17276 9163
rect 17224 9120 17276 9129
rect 18328 9120 18380 9172
rect 20444 9163 20496 9172
rect 20444 9129 20453 9163
rect 20453 9129 20487 9163
rect 20487 9129 20496 9163
rect 20444 9120 20496 9129
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 10784 8984 10836 9036
rect 16396 8984 16448 9036
rect 17868 9027 17920 9036
rect 17868 8993 17877 9027
rect 17877 8993 17911 9027
rect 17911 8993 17920 9027
rect 17868 8984 17920 8993
rect 13268 8916 13320 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 15568 8916 15620 8968
rect 16948 8916 17000 8968
rect 21364 8959 21416 8968
rect 11888 8848 11940 8900
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 15568 8780 15620 8832
rect 17500 8780 17552 8832
rect 18328 8823 18380 8832
rect 18328 8789 18337 8823
rect 18337 8789 18371 8823
rect 18371 8789 18380 8823
rect 18328 8780 18380 8789
rect 18972 8780 19024 8832
rect 20996 8823 21048 8832
rect 20996 8789 21005 8823
rect 21005 8789 21039 8823
rect 21039 8789 21048 8823
rect 20996 8780 21048 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 5816 8576 5868 8628
rect 11888 8576 11940 8628
rect 13268 8619 13320 8628
rect 7840 8508 7892 8560
rect 10692 8508 10744 8560
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 9588 8440 9640 8492
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 11152 8508 11204 8560
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 15108 8619 15160 8628
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 18512 8576 18564 8628
rect 20076 8576 20128 8628
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 15936 8483 15988 8492
rect 15936 8449 15945 8483
rect 15945 8449 15979 8483
rect 15979 8449 15988 8483
rect 15936 8440 15988 8449
rect 18052 8440 18104 8492
rect 18880 8440 18932 8492
rect 10416 8372 10468 8381
rect 11152 8372 11204 8424
rect 12716 8415 12768 8424
rect 8116 8347 8168 8356
rect 8116 8313 8125 8347
rect 8125 8313 8159 8347
rect 8159 8313 8168 8347
rect 8116 8304 8168 8313
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 14372 8372 14424 8424
rect 14648 8415 14700 8424
rect 12992 8304 13044 8356
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 14648 8372 14700 8381
rect 17040 8347 17092 8356
rect 17040 8313 17049 8347
rect 17049 8313 17083 8347
rect 17083 8313 17092 8347
rect 17040 8304 17092 8313
rect 7840 8279 7892 8288
rect 7840 8245 7849 8279
rect 7849 8245 7883 8279
rect 7883 8245 7892 8279
rect 7840 8236 7892 8245
rect 9404 8236 9456 8288
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 20720 8508 20772 8560
rect 19524 8304 19576 8356
rect 21180 8304 21232 8356
rect 21364 8347 21416 8356
rect 21364 8313 21373 8347
rect 21373 8313 21407 8347
rect 21407 8313 21416 8347
rect 21364 8304 21416 8313
rect 17960 8236 18012 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 9128 8032 9180 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 14372 8032 14424 8084
rect 18880 8032 18932 8084
rect 10416 7964 10468 8016
rect 16948 7964 17000 8016
rect 18512 8007 18564 8016
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 11888 7896 11940 7948
rect 18512 7973 18521 8007
rect 18521 7973 18555 8007
rect 18555 7973 18564 8007
rect 18512 7964 18564 7973
rect 17684 7939 17736 7948
rect 17684 7905 17693 7939
rect 17693 7905 17727 7939
rect 17727 7905 17736 7939
rect 17684 7896 17736 7905
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 13820 7828 13872 7880
rect 17960 7760 18012 7812
rect 8208 7692 8260 7744
rect 14924 7692 14976 7744
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 9588 7488 9640 7540
rect 13636 7488 13688 7540
rect 18420 7488 18472 7540
rect 20352 7488 20404 7540
rect 8300 7420 8352 7472
rect 9404 7420 9456 7472
rect 9496 7420 9548 7472
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 20536 7420 20588 7472
rect 7288 7284 7340 7336
rect 21088 7395 21140 7404
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18052 7284 18104 7336
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 17132 7216 17184 7268
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 10692 6944 10744 6996
rect 15476 6944 15528 6996
rect 1584 6808 1636 6860
rect 9588 6876 9640 6928
rect 11152 6876 11204 6928
rect 9404 6740 9456 6792
rect 10600 6740 10652 6792
rect 11796 6808 11848 6860
rect 17408 6808 17460 6860
rect 11520 6740 11572 6792
rect 13176 6740 13228 6792
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 14648 6672 14700 6724
rect 21272 6740 21324 6792
rect 9312 6604 9364 6613
rect 10784 6604 10836 6656
rect 12532 6604 12584 6656
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 15936 6604 15988 6656
rect 19616 6604 19668 6656
rect 19892 6647 19944 6656
rect 19892 6613 19901 6647
rect 19901 6613 19935 6647
rect 19935 6613 19944 6647
rect 19892 6604 19944 6613
rect 20444 6647 20496 6656
rect 20444 6613 20453 6647
rect 20453 6613 20487 6647
rect 20487 6613 20496 6647
rect 20444 6604 20496 6613
rect 20812 6604 20864 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 9312 6400 9364 6452
rect 9404 6400 9456 6452
rect 10508 6400 10560 6452
rect 10784 6443 10836 6452
rect 10784 6409 10793 6443
rect 10793 6409 10827 6443
rect 10827 6409 10836 6443
rect 10784 6400 10836 6409
rect 13820 6400 13872 6452
rect 15384 6400 15436 6452
rect 17316 6400 17368 6452
rect 21088 6400 21140 6452
rect 16396 6332 16448 6384
rect 8484 6264 8536 6316
rect 9496 6264 9548 6316
rect 11152 6264 11204 6316
rect 11704 6264 11756 6316
rect 11980 6264 12032 6316
rect 11060 6239 11112 6248
rect 9588 6128 9640 6180
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 12532 6196 12584 6248
rect 12440 6128 12492 6180
rect 13636 6128 13688 6180
rect 19064 6264 19116 6316
rect 16028 6196 16080 6248
rect 15384 6128 15436 6180
rect 8208 6060 8260 6112
rect 11980 6060 12032 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 9496 5856 9548 5908
rect 11704 5763 11756 5772
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 13084 5720 13136 5772
rect 12256 5652 12308 5704
rect 18052 5720 18104 5772
rect 4068 5584 4120 5636
rect 15016 5584 15068 5636
rect 9496 5516 9548 5568
rect 12440 5516 12492 5568
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 21272 5559 21324 5568
rect 21272 5525 21281 5559
rect 21281 5525 21315 5559
rect 21315 5525 21324 5559
rect 21272 5516 21324 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 1492 5312 1544 5364
rect 12624 5312 12676 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 15292 5312 15344 5321
rect 15568 5312 15620 5364
rect 18144 5312 18196 5364
rect 11060 5176 11112 5228
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 9496 5108 9548 5160
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 15752 5151 15804 5160
rect 13636 5108 13688 5117
rect 15752 5117 15761 5151
rect 15761 5117 15795 5151
rect 15795 5117 15804 5151
rect 15752 5108 15804 5117
rect 16028 5108 16080 5160
rect 18696 5040 18748 5092
rect 9220 4972 9272 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 12256 5015 12308 5024
rect 12256 4981 12265 5015
rect 12265 4981 12299 5015
rect 12299 4981 12308 5015
rect 12256 4972 12308 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 13176 4811 13228 4820
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 9496 4632 9548 4684
rect 10692 4632 10744 4684
rect 12256 4632 12308 4684
rect 13176 4777 13185 4811
rect 13185 4777 13219 4811
rect 13219 4777 13228 4811
rect 13176 4768 13228 4777
rect 14740 4564 14792 4616
rect 8392 4496 8444 4548
rect 11520 4496 11572 4548
rect 11888 4496 11940 4548
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 12072 4428 12124 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 9312 4224 9364 4276
rect 10048 4224 10100 4276
rect 10784 4224 10836 4276
rect 12072 4267 12124 4276
rect 9496 4156 9548 4208
rect 1400 4020 1452 4072
rect 8668 4020 8720 4072
rect 9496 4020 9548 4072
rect 10600 4088 10652 4140
rect 11060 4156 11112 4208
rect 12072 4233 12081 4267
rect 12081 4233 12115 4267
rect 12115 4233 12124 4267
rect 12072 4224 12124 4233
rect 12532 4224 12584 4276
rect 17960 4224 18012 4276
rect 10600 3952 10652 4004
rect 11152 3995 11204 4004
rect 11152 3961 11161 3995
rect 11161 3961 11195 3995
rect 11195 3961 11204 3995
rect 11152 3952 11204 3961
rect 11888 3952 11940 4004
rect 16396 4088 16448 4140
rect 18052 4088 18104 4140
rect 17960 4020 18012 4072
rect 13820 3995 13872 4004
rect 13820 3961 13829 3995
rect 13829 3961 13863 3995
rect 13863 3961 13872 3995
rect 13820 3952 13872 3961
rect 14556 3952 14608 4004
rect 18972 3952 19024 4004
rect 15476 3884 15528 3936
rect 17592 3884 17644 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 9496 3680 9548 3732
rect 10048 3680 10100 3732
rect 10600 3723 10652 3732
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 11060 3680 11112 3732
rect 15660 3680 15712 3732
rect 15752 3680 15804 3732
rect 17592 3680 17644 3732
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 17776 3544 17828 3596
rect 17040 3476 17092 3528
rect 14556 3340 14608 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 15568 3383 15620 3392
rect 14648 3340 14700 3349
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 15660 3383 15712 3392
rect 15660 3349 15669 3383
rect 15669 3349 15703 3383
rect 15703 3349 15712 3383
rect 15660 3340 15712 3349
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 12164 3136 12216 3188
rect 15568 3136 15620 3188
rect 14648 3000 14700 3052
rect 17960 3000 18012 3052
rect 15660 2796 15712 2848
rect 19064 2796 19116 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 15384 2592 15436 2644
rect 19156 2592 19208 2644
rect 12440 2524 12492 2576
rect 19248 2524 19300 2576
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
<< metal2 >>
rect 386 22200 442 23000
rect 938 22200 994 23000
rect 1490 22200 1546 23000
rect 1596 22222 1992 22250
rect 400 18426 428 22200
rect 952 19242 980 22200
rect 1400 19440 1452 19446
rect 1400 19382 1452 19388
rect 940 19236 992 19242
rect 940 19178 992 19184
rect 388 18420 440 18426
rect 388 18362 440 18368
rect 1412 4078 1440 19382
rect 1504 5370 1532 22200
rect 1596 6866 1624 22222
rect 1964 22114 1992 22222
rect 2042 22200 2098 23000
rect 2594 22200 2650 23000
rect 3146 22200 3202 23000
rect 3698 22200 3754 23000
rect 3804 22222 4016 22250
rect 2056 22114 2084 22200
rect 1964 22086 2084 22114
rect 2608 19446 2636 22200
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 3160 18970 3188 22200
rect 3712 22114 3740 22200
rect 3804 22114 3832 22222
rect 3712 22086 3832 22114
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3882 19816 3938 19825
rect 3882 19751 3938 19760
rect 3896 19514 3924 19751
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3988 19310 4016 22222
rect 4250 22200 4306 23000
rect 4802 22200 4858 23000
rect 5354 22200 5410 23000
rect 5906 22200 5962 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7116 22222 7512 22250
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4264 19802 4292 22200
rect 4712 19848 4764 19854
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2424 16454 2452 18702
rect 4172 18698 4200 19790
rect 4264 19774 4476 19802
rect 4712 19790 4764 19796
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3884 17740 3936 17746
rect 3884 17682 3936 17688
rect 3896 17241 3924 17682
rect 3882 17232 3938 17241
rect 3882 17167 3938 17176
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 4264 14074 4292 19382
rect 4356 19174 4384 19654
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17338 4384 17478
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 4448 13530 4476 19774
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4540 18358 4568 19314
rect 4528 18352 4580 18358
rect 4528 18294 4580 18300
rect 4724 17882 4752 19790
rect 4816 19446 4844 22200
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 5368 19334 5396 22200
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5736 20058 5764 20266
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5920 19394 5948 22200
rect 6472 20890 6500 22200
rect 6472 20862 6592 20890
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 5736 19366 5948 19394
rect 5368 19306 5580 19334
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4816 17338 4844 18226
rect 4908 18154 4936 18634
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4540 14822 4568 16594
rect 5184 15162 5212 18702
rect 5552 16454 5580 19306
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5644 17338 5672 17682
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5552 16250 5580 16390
rect 5736 16250 5764 19366
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 5644 14482 5672 14962
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 5736 9042 5764 9386
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5828 8634 5856 19178
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6472 17898 6500 18362
rect 6564 18086 6592 20862
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 5908 17876 5960 17882
rect 6472 17870 6592 17898
rect 5908 17818 5960 17824
rect 5920 17134 5948 17818
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 6012 16658 6040 17614
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6012 16182 6040 16458
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6564 9518 6592 17870
rect 6656 9654 6684 19246
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 16794 6868 18158
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 17202 6960 18022
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16794 6960 17138
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7024 16574 7052 22200
rect 6932 16546 7052 16574
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6748 13258 6776 16118
rect 6840 15162 6868 16390
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6748 11898 6776 12038
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6840 11694 6868 12038
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4080 5642 4108 5743
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 6932 5273 6960 16546
rect 7116 15094 7144 22222
rect 7484 22114 7512 22222
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10520 22222 10824 22250
rect 7576 22114 7604 22200
rect 7484 22086 7604 22114
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7300 19446 7328 20470
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7208 16454 7236 17546
rect 7300 16522 7328 18022
rect 7288 16516 7340 16522
rect 7288 16458 7340 16464
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7300 13326 7328 13466
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 11830 7052 13126
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7116 10130 7144 10610
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7300 8430 7328 11494
rect 7392 11354 7420 18906
rect 7576 12986 7604 19314
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7760 18290 7788 18634
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7852 17270 7880 18566
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7668 14822 7696 14962
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7392 10742 7420 11290
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7668 9586 7696 14758
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7300 7342 7328 8366
rect 7760 7546 7788 13466
rect 7852 8566 7880 16390
rect 8128 15162 8156 22200
rect 8680 18766 8708 22200
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9140 18834 9168 19858
rect 9232 19394 9260 22200
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 19922 9352 20334
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9232 19366 9444 19394
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8220 14634 8248 18566
rect 8680 18426 8708 18702
rect 9048 18426 9076 18702
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8496 16574 8524 17546
rect 8404 16546 8524 16574
rect 8404 16114 8432 16546
rect 8680 16454 8708 18226
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9232 16794 9260 17682
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8404 15910 8432 16050
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8036 14606 8248 14634
rect 8036 13530 8064 14606
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 14074 8156 14214
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8220 10810 8248 14418
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8220 10470 8248 10746
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8128 10062 8156 10406
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8220 9874 8248 10406
rect 8128 9846 8248 9874
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 8128 8362 8156 9846
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 7954 7880 8230
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 8128 6644 8156 8298
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7546 8248 7686
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7478 8340 13194
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 6656 8260 6662
rect 8128 6616 8208 6644
rect 8208 6598 8260 6604
rect 8220 6118 8248 6598
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 8404 4554 8432 15846
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9324 14074 9352 18158
rect 9416 14074 9444 19366
rect 9784 19310 9812 22200
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9508 16658 9536 18022
rect 10244 17882 10272 19654
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 9588 17808 9640 17814
rect 9640 17756 9720 17762
rect 9588 17750 9720 17756
rect 9600 17734 9720 17750
rect 10336 17746 10364 22200
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 9692 17542 9720 17734
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9600 17218 9628 17478
rect 10428 17338 10456 19314
rect 10520 17542 10548 22222
rect 10796 22114 10824 22222
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 11532 22222 11928 22250
rect 10888 22114 10916 22200
rect 10796 22086 10916 22114
rect 11440 22114 11468 22200
rect 11532 22114 11560 22222
rect 11440 22086 11560 22114
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 9600 17190 9720 17218
rect 9692 17066 9720 17190
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14550 9720 14758
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9416 10062 9444 10542
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9722 9352 9862
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8496 6322 8524 7346
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 8680 4078 8708 9522
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 9140 8090 9168 8366
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9416 7886 9444 8230
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9508 7478 9536 14214
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 13297 9628 13670
rect 9784 13530 9812 17070
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16250 10088 16390
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9968 14414 9996 15030
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9586 13288 9642 13297
rect 9586 13223 9642 13232
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 8498 9628 12582
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9416 6798 9444 7414
rect 9600 6934 9628 7482
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6458 9352 6598
rect 9416 6458 9444 6734
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9508 5914 9536 6258
rect 9600 6186 9628 6870
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9508 5574 9536 5850
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9232 4690 9260 4966
rect 9508 4690 9536 5102
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9508 4214 9536 4626
rect 10060 4282 10088 13806
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12986 10456 13126
rect 10520 12986 10548 14214
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10152 11354 10180 12174
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10612 10130 10640 20402
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18358 10732 18566
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10704 17610 10732 18294
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10704 9178 10732 14010
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10796 9042 10824 19314
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10888 13530 10916 19246
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11072 18358 11100 18634
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10980 16658 11008 18226
rect 11164 17066 11192 18634
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10888 13326 10916 13466
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11164 11626 11192 12854
rect 11256 12306 11284 19790
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11716 19446 11744 19790
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11900 19394 11928 22222
rect 11978 22200 12034 23000
rect 12530 22200 12586 23000
rect 13082 22200 13138 23000
rect 13188 22222 13584 22250
rect 11992 20058 12020 22200
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 11520 19372 11572 19378
rect 11900 19366 12112 19394
rect 11520 19314 11572 19320
rect 11532 19174 11560 19314
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11716 18154 11744 18566
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11624 16658 11652 17138
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11808 16574 11836 17138
rect 11808 16546 11928 16574
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11716 14618 11744 16458
rect 11900 15366 11928 16546
rect 11992 16250 12020 18634
rect 12084 16574 12112 19366
rect 12268 17921 12296 19858
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12452 18426 12480 18702
rect 12544 18426 12572 22200
rect 13096 20602 13124 22200
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13188 19530 13216 22222
rect 13556 22114 13584 22222
rect 13634 22200 13690 23000
rect 13832 22222 14136 22250
rect 13648 22114 13676 22200
rect 13556 22086 13676 22114
rect 13832 19530 13860 22222
rect 14108 22114 14136 22222
rect 14186 22200 14242 23000
rect 14738 22200 14794 23000
rect 14844 22222 15148 22250
rect 14200 22114 14228 22200
rect 14108 22086 14228 22114
rect 14752 22114 14780 22200
rect 14844 22114 14872 22222
rect 14752 22086 14872 22114
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 12636 19502 13216 19530
rect 13740 19514 13860 19530
rect 13728 19508 13860 19514
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12348 18080 12400 18086
rect 12346 18048 12348 18057
rect 12400 18048 12402 18057
rect 12346 17983 12402 17992
rect 12254 17912 12310 17921
rect 12254 17847 12310 17856
rect 12452 17678 12480 18362
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12452 17270 12480 17614
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12360 16794 12388 17138
rect 12636 16810 12664 19502
rect 13780 19502 13860 19508
rect 13728 19450 13780 19456
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12452 16782 12664 16810
rect 12084 16546 12204 16574
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16250 12112 16390
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13462 11652 13670
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10606 11100 10950
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10428 8022 10456 8366
rect 10704 8090 10732 8502
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10520 6458 10548 7346
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 9508 3738 9536 4014
rect 10060 3738 10088 4218
rect 10612 4146 10640 6734
rect 10704 4690 10732 6938
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6458 10824 6598
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11072 6254 11100 10542
rect 11164 8566 11192 11562
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11716 9926 11744 13806
rect 11900 13802 11928 15302
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11256 9518 11284 9862
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11164 6934 11192 8366
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11532 6798 11560 7278
rect 11808 6866 11836 11018
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8634 11928 8842
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 7954 11928 8434
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10796 4282 10824 4422
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 11072 4214 11100 5170
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10612 3738 10640 3946
rect 11072 3738 11100 4150
rect 11164 4010 11192 6258
rect 11716 5778 11744 6258
rect 11992 6118 12020 6258
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4554 11560 4966
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11900 4010 11928 4490
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4282 12112 4422
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 12176 3194 12204 16546
rect 12452 14414 12480 16782
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12360 11082 12388 12378
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12268 9586 12296 9998
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12360 9178 12388 9386
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 6186 12480 13194
rect 12544 12850 12572 16390
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12728 12434 12756 18362
rect 12912 16454 12940 19382
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13280 19174 13308 19246
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18766 13768 19110
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13188 17882 13216 18634
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13648 18290 13676 18566
rect 13740 18426 13768 18702
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13740 18290 13768 18362
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13740 17882 13768 18226
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 13820 18080 13872 18086
rect 13818 18048 13820 18057
rect 13872 18048 13874 18057
rect 13818 17983 13874 17992
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13818 17912 13874 17921
rect 13945 17915 14253 17924
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13728 17876 13780 17882
rect 13818 17847 13874 17856
rect 13728 17818 13780 17824
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 17066 13124 17614
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 13004 16114 13032 16934
rect 13188 16182 13216 17818
rect 13832 17762 13860 17847
rect 14292 17762 14320 18090
rect 13832 17734 14320 17762
rect 13832 16454 13860 17734
rect 14384 17202 14412 19314
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13176 16176 13228 16182
rect 13176 16118 13228 16124
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 14822 13032 16050
rect 13464 15910 13492 16390
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13464 15502 13492 15846
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 13190 13124 14282
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13188 12434 13216 15370
rect 13464 15366 13492 15438
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14278 13492 15302
rect 14292 14822 14320 15506
rect 14384 14958 14412 17138
rect 15120 16574 15148 22222
rect 15290 22200 15346 23000
rect 15396 22222 15608 22250
rect 15304 22114 15332 22200
rect 15396 22114 15424 22222
rect 15304 22086 15424 22114
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 18358 15240 19790
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15212 16590 15240 16934
rect 15028 16546 15148 16574
rect 15200 16584 15252 16590
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13464 14006 13492 14214
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13464 13870 13492 13942
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13464 13530 13492 13806
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13464 13326 13492 13466
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13372 12434 13400 13126
rect 13464 12986 13492 13262
rect 13740 13258 13768 14214
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 12636 12406 12756 12434
rect 13004 12406 13216 12434
rect 13280 12406 13400 12434
rect 12636 6905 12664 12406
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12728 10266 12756 12106
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11558 12848 11834
rect 13004 11558 13032 12406
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12912 11257 12940 11290
rect 12898 11248 12954 11257
rect 12898 11183 12954 11192
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10810 12940 10950
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12912 10062 12940 10746
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 8430 12756 9318
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 13004 8362 13032 11494
rect 13280 11234 13308 12406
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11354 13400 11562
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13096 11206 13308 11234
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12622 6896 12678 6905
rect 12622 6831 12678 6840
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6254 12572 6598
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12544 6118 12572 6190
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12268 5710 12296 6054
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12268 4690 12296 4966
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 12452 2582 12480 5510
rect 12544 4282 12572 6054
rect 13096 5778 13124 11206
rect 13464 11150 13492 12922
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13280 10810 13308 11086
rect 13556 11014 13584 13126
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13280 10266 13308 10746
rect 13648 10470 13676 11698
rect 13832 11082 13860 12582
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 14292 12102 14320 14758
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8634 13308 8910
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13648 7546 13676 10406
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 7886 13860 9590
rect 14476 9450 14504 15846
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12434 14872 13126
rect 15028 12434 15056 16546
rect 15200 16526 15252 16532
rect 15304 16522 15332 18022
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15212 14890 15240 16390
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15212 14346 15240 14826
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 14752 12406 14872 12434
rect 14936 12406 15056 12434
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14200 8945 14228 9114
rect 14568 8974 14596 11766
rect 14752 10674 14780 12406
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14556 8968 14608 8974
rect 14186 8936 14242 8945
rect 14556 8910 14608 8916
rect 14186 8871 14242 8880
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14384 8090 14412 8366
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5370 12664 5510
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12714 5264 12770 5273
rect 12714 5199 12716 5208
rect 12768 5199 12770 5208
rect 12716 5170 12768 5176
rect 13188 4826 13216 6734
rect 14660 6730 14688 8366
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 5166 13676 6122
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 13832 4010 13860 6394
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 14752 4622 14780 10610
rect 14936 7750 14964 12406
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15212 11830 15240 12106
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 11082 15056 11494
rect 15304 11257 15332 12106
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15028 10674 15056 11018
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15028 5642 15056 9862
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15120 8634 15148 9522
rect 15212 9160 15240 10950
rect 15304 10266 15332 11183
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15292 9172 15344 9178
rect 15212 9132 15292 9160
rect 15292 9114 15344 9120
rect 15396 9081 15424 19382
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15488 16998 15516 18634
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15488 16794 15516 16934
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15580 15144 15608 22222
rect 15842 22200 15898 23000
rect 16394 22200 16450 23000
rect 16946 22200 17002 23000
rect 17498 22200 17554 23000
rect 18050 22200 18106 23000
rect 18602 22200 18658 23000
rect 19154 22200 19210 23000
rect 19706 22200 19762 23000
rect 20258 22200 20314 23000
rect 20810 22200 20866 23000
rect 21362 22200 21418 23000
rect 21560 22222 21864 22250
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15764 16590 15792 17206
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15580 15116 15792 15144
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15488 14074 15516 14282
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 11286 15516 12718
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15382 9072 15438 9081
rect 15382 9007 15438 9016
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15488 7002 15516 11222
rect 15580 10470 15608 13194
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15672 9450 15700 12582
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15568 8968 15620 8974
rect 15566 8936 15568 8945
rect 15764 8945 15792 15116
rect 15856 9489 15884 22200
rect 16408 19446 16436 22200
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16960 19394 16988 22200
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17328 19854 17356 20334
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 16960 19366 17080 19394
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16316 18630 16344 18906
rect 16960 18630 16988 19246
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16224 14618 16252 14962
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16224 13870 16252 14554
rect 16408 14550 16436 15030
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 13530 16252 13806
rect 16408 13802 16436 14486
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12442 16068 13126
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 16960 12238 16988 18362
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16028 12096 16080 12102
rect 17052 12050 17080 19366
rect 17144 18698 17172 19790
rect 17512 18850 17540 22200
rect 17866 21040 17922 21049
rect 17866 20975 17922 20984
rect 17880 20058 17908 20975
rect 17958 20496 18014 20505
rect 17958 20431 18014 20440
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17972 19990 18000 20431
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17420 18822 17540 18850
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17328 17678 17356 18566
rect 17420 18426 17448 18822
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17512 18154 17540 18634
rect 17500 18148 17552 18154
rect 17500 18090 17552 18096
rect 17696 17785 17724 19654
rect 17682 17776 17738 17785
rect 17682 17711 17738 17720
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17604 16250 17632 16458
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17316 14408 17368 14414
rect 17236 14356 17316 14362
rect 17236 14350 17368 14356
rect 17236 14334 17356 14350
rect 17236 12434 17264 14334
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17604 13326 17632 13670
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17696 12714 17724 15302
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17696 12594 17724 12650
rect 16028 12038 16080 12044
rect 15842 9480 15898 9489
rect 15842 9415 15898 9424
rect 15620 8936 15622 8945
rect 15566 8871 15622 8880
rect 15750 8936 15806 8945
rect 15750 8871 15806 8880
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15304 5370 15332 6598
rect 15396 6458 15424 6598
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14568 3602 14596 3946
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14568 3398 14596 3538
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14660 3058 14688 3334
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 15396 2650 15424 6122
rect 15580 5370 15608 8774
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15948 6662 15976 8434
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16040 6254 16068 12038
rect 16960 12022 17080 12050
rect 17144 12406 17264 12434
rect 17604 12566 17724 12594
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10062 16528 10406
rect 16488 10056 16540 10062
rect 16408 10004 16488 10010
rect 16408 9998 16540 10004
rect 16408 9982 16528 9998
rect 16408 9042 16436 9982
rect 16868 9926 16896 10610
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16960 9058 16988 12022
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17052 11150 17080 11834
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17144 9382 17172 12406
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 9874 17264 12174
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10742 17356 11086
rect 17420 10810 17448 11494
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17328 10130 17356 10678
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17236 9846 17356 9874
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17236 9178 17264 9658
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 16396 9036 16448 9042
rect 16960 9030 17172 9058
rect 16396 8978 16448 8984
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 8022 16988 8910
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15488 3602 15516 3878
rect 15672 3738 15700 5170
rect 16040 5166 16068 6190
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 15764 3738 15792 5102
rect 16408 4146 16436 6326
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 17052 3534 17080 8298
rect 17144 7274 17172 9030
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17328 6458 17356 9846
rect 17420 6866 17448 10746
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17512 5545 17540 8774
rect 17498 5536 17554 5545
rect 17498 5471 17554 5480
rect 17604 3942 17632 12566
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17696 7954 17724 11290
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17604 3738 17632 3878
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17788 3602 17816 19790
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17880 18766 17908 19382
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17880 18222 17908 18702
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17880 17882 17908 18158
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17880 17338 17908 17818
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17880 16658 17908 17274
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 16250 17908 16594
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17880 15502 17908 16186
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17880 15162 17908 15438
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 18064 13530 18092 22200
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 18737 18184 20198
rect 18616 20058 18644 22200
rect 19168 20346 19196 22200
rect 18984 20318 19196 20346
rect 19616 20324 19668 20330
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18800 19854 18828 20198
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18142 18728 18198 18737
rect 18142 18663 18198 18672
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18156 17610 18184 18226
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17958 13424 18014 13433
rect 18156 13410 18184 15370
rect 17958 13359 18014 13368
rect 18064 13382 18184 13410
rect 17972 12646 18000 13359
rect 18064 13258 18092 13382
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18064 12458 18092 13194
rect 17972 12430 18092 12458
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17880 9042 17908 11766
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17972 8294 18000 12430
rect 18248 11257 18276 19790
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18432 17241 18460 19722
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18418 17232 18474 17241
rect 18418 17167 18474 17176
rect 18326 15600 18382 15609
rect 18326 15535 18382 15544
rect 18234 11248 18290 11257
rect 18234 11183 18290 11192
rect 18340 9178 18368 15535
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18432 12986 18460 13262
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18524 12753 18552 19314
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18616 18873 18644 19110
rect 18602 18864 18658 18873
rect 18602 18799 18658 18808
rect 18708 18290 18736 19110
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18694 14920 18750 14929
rect 18694 14855 18750 14864
rect 18510 12744 18566 12753
rect 18510 12679 18566 12688
rect 18708 12434 18736 14855
rect 18786 13152 18842 13161
rect 18786 13087 18842 13096
rect 18524 12406 18736 12434
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18432 12102 18460 12174
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11762 18460 12038
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18524 10690 18552 12406
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11830 18736 12038
rect 18696 11824 18748 11830
rect 18696 11766 18748 11772
rect 18708 11694 18736 11766
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18708 11150 18736 11630
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18432 10662 18552 10690
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 18064 7954 18092 8434
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17972 7342 18000 7754
rect 17960 7336 18012 7342
rect 17958 7304 17960 7313
rect 18052 7336 18104 7342
rect 18012 7304 18014 7313
rect 18052 7278 18104 7284
rect 17958 7239 18014 7248
rect 18064 5778 18092 7278
rect 18340 6361 18368 8774
rect 18432 7546 18460 10662
rect 18800 10554 18828 13087
rect 18892 12889 18920 20198
rect 18984 18426 19012 20318
rect 19616 20266 19668 20272
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19246 19952 19302 19961
rect 19246 19887 19248 19896
rect 19300 19887 19302 19896
rect 19248 19858 19300 19864
rect 19524 19848 19576 19854
rect 19628 19825 19656 20266
rect 19720 19990 19748 22200
rect 20272 20058 20300 22200
rect 20626 21448 20682 21457
rect 20626 21383 20682 21392
rect 20640 20602 20668 21383
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 19708 19984 19760 19990
rect 19708 19926 19760 19932
rect 20640 19854 20668 20538
rect 20824 19990 20852 22200
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20260 19848 20312 19854
rect 19524 19790 19576 19796
rect 19614 19816 19670 19825
rect 19536 19242 19564 19790
rect 20260 19790 20312 19796
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 19614 19751 19670 19760
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 20272 19174 20300 19790
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 19076 18766 19104 19110
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19536 18086 19564 18634
rect 19524 18080 19576 18086
rect 19522 18048 19524 18057
rect 19576 18048 19578 18057
rect 19143 17980 19451 17989
rect 19522 17983 19578 17992
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17202 19748 17478
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 18970 16144 19026 16153
rect 18970 16079 19026 16088
rect 18878 12880 18934 12889
rect 18878 12815 18934 12824
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18524 10526 18828 10554
rect 18524 8634 18552 10526
rect 18892 10282 18920 12582
rect 18708 10254 18920 10282
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18524 8022 18552 8366
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18326 6352 18382 6361
rect 18326 6287 18382 6296
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 17958 4720 18014 4729
rect 17958 4655 18014 4664
rect 17972 4282 18000 4655
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 18156 4185 18184 5306
rect 18708 5098 18736 10254
rect 18878 10160 18934 10169
rect 18878 10095 18934 10104
rect 18892 8498 18920 10095
rect 18984 8838 19012 16079
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19076 15473 19104 15846
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19062 15464 19118 15473
rect 19062 15399 19118 15408
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19536 14822 19564 15370
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19248 14612 19300 14618
rect 19300 14572 19380 14600
rect 19248 14554 19300 14560
rect 19352 13870 19380 14572
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19340 13184 19392 13190
rect 19260 13132 19340 13138
rect 19260 13126 19392 13132
rect 19260 13110 19380 13126
rect 19260 12646 19288 13110
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19076 11218 19104 11834
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19168 10810 19196 11018
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19062 9616 19118 9625
rect 19062 9551 19118 9560
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18892 8090 18920 8434
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 19076 6322 19104 9551
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19536 8362 19564 14758
rect 19614 13968 19670 13977
rect 19614 13903 19670 13912
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19628 6662 19656 13903
rect 19720 13734 19748 17138
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19890 14512 19946 14521
rect 19890 14447 19946 14456
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11762 19840 12038
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19904 9450 19932 14447
rect 19996 14414 20024 15846
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 12238 20024 12582
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 20088 8634 20116 13806
rect 20272 12209 20300 19110
rect 20350 18184 20406 18193
rect 20350 18119 20406 18128
rect 20258 12200 20314 12209
rect 20258 12135 20314 12144
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20364 7546 20392 18119
rect 20456 11665 20484 19178
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20916 17678 20944 18294
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20902 16960 20958 16969
rect 20902 16895 20958 16904
rect 20916 16794 20944 16895
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 21008 16574 21036 19382
rect 21192 19378 21220 20198
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21284 19174 21312 19858
rect 21376 19514 21404 22200
rect 21560 20602 21588 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22466 22200 22522 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 22480 19446 22508 22200
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18766 21312 19110
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18358 21220 18566
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21284 18086 21312 18702
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21284 17678 21312 18022
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21284 16998 21312 17614
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21284 16658 21312 16934
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 20626 16552 20682 16561
rect 20626 16487 20682 16496
rect 20916 16546 21036 16574
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20442 11656 20498 11665
rect 20442 11591 20498 11600
rect 20548 11354 20576 16050
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20442 9480 20498 9489
rect 20442 9415 20498 9424
rect 20456 9178 20484 9415
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20442 8936 20498 8945
rect 20442 8871 20498 8880
rect 20456 8634 20484 8871
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20548 7478 20576 9522
rect 20640 9450 20668 16487
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20732 14278 20760 15030
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20732 8566 20760 14214
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20824 13394 20852 14010
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20824 12918 20852 13330
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20916 12434 20944 16546
rect 21284 16114 21312 16594
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21284 15706 21312 16050
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21284 15026 21312 15642
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 14618 21312 14962
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21284 14074 21312 14554
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21192 13326 21220 13670
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20824 12406 20944 12434
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 19890 6896 19946 6905
rect 19890 6831 19946 6840
rect 19904 6662 19932 6831
rect 20824 6662 20852 12406
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 11354 20944 11698
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20916 10810 20944 11290
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21192 10033 21220 13262
rect 21272 12912 21324 12918
rect 21272 12854 21324 12860
rect 21284 12238 21312 12854
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11762 21312 12174
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21468 10713 21496 18226
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21454 10704 21510 10713
rect 21272 10668 21324 10674
rect 21454 10639 21510 10648
rect 21272 10610 21324 10616
rect 21284 10266 21312 10610
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21178 10024 21234 10033
rect 21178 9959 21234 9968
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21086 9208 21142 9217
rect 21086 9143 21142 9152
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 8401 21036 8774
rect 20994 8392 21050 8401
rect 20994 8327 21050 8336
rect 21100 7410 21128 9143
rect 21192 9081 21220 9318
rect 21178 9072 21234 9081
rect 21178 9007 21234 9016
rect 21376 8974 21404 9522
rect 21364 8968 21416 8974
rect 21362 8936 21364 8945
rect 21416 8936 21418 8945
rect 21362 8871 21418 8880
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 20456 5953 20484 6598
rect 21100 6458 21128 7346
rect 21192 6769 21220 8298
rect 21376 7993 21404 8298
rect 21362 7984 21418 7993
rect 21362 7919 21418 7928
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 7449 21312 7686
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21270 7440 21326 7449
rect 21270 7375 21326 7384
rect 21272 6792 21324 6798
rect 21178 6760 21234 6769
rect 21272 6734 21324 6740
rect 21178 6695 21234 6704
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20442 5944 20498 5953
rect 20442 5879 20498 5888
rect 21284 5574 21312 6734
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21284 5137 21312 5510
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21270 5128 21326 5137
rect 18696 5092 18748 5098
rect 21270 5063 21326 5072
rect 18696 5034 18748 5040
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 18142 4176 18198 4185
rect 18052 4140 18104 4146
rect 18142 4111 18198 4120
rect 18052 4082 18104 4088
rect 17960 4072 18012 4078
rect 17958 4040 17960 4049
rect 18012 4040 18014 4049
rect 17958 3975 18014 3984
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17040 3528 17092 3534
rect 18064 3505 18092 4082
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 17040 3470 17092 3476
rect 18050 3496 18106 3505
rect 18050 3431 18106 3440
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15580 3194 15608 3334
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15672 2854 15700 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 17958 3088 18014 3097
rect 17958 3023 17960 3032
rect 18012 3023 18014 3032
rect 17960 2994 18012 3000
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 18984 2417 19012 3946
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18970 2408 19026 2417
rect 18970 2343 19026 2352
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 19076 1465 19104 2790
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19168 1873 19196 2586
rect 19248 2576 19300 2582
rect 19246 2544 19248 2553
rect 19300 2544 19302 2553
rect 19246 2479 19302 2488
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 19154 1864 19210 1873
rect 19154 1799 19210 1808
rect 19062 1456 19118 1465
rect 19062 1391 19118 1400
<< via2 >>
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3882 19760 3938 19816
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3882 17176 3938 17232
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 4066 5752 4122 5808
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 6918 5208 6974 5264
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9586 13232 9642 13288
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12346 18028 12348 18048
rect 12348 18028 12400 18048
rect 12400 18028 12402 18048
rect 12346 17992 12402 18028
rect 12254 17856 12310 17912
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13818 18028 13820 18048
rect 13820 18028 13872 18048
rect 13872 18028 13874 18048
rect 13818 17992 13874 18028
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13818 17856 13874 17912
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 12898 11192 12954 11248
rect 12622 6840 12678 6896
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14186 8880 14242 8936
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 12714 5228 12770 5264
rect 12714 5208 12716 5228
rect 12716 5208 12768 5228
rect 12768 5208 12770 5228
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 15290 11192 15346 11248
rect 15382 9016 15438 9072
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 17866 20984 17922 21040
rect 17958 20440 18014 20496
rect 17682 17720 17738 17776
rect 15842 9424 15898 9480
rect 15566 8916 15568 8936
rect 15568 8916 15620 8936
rect 15620 8916 15622 8936
rect 15566 8880 15622 8916
rect 15750 8880 15806 8936
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 17498 5480 17554 5536
rect 18142 18672 18198 18728
rect 17958 13368 18014 13424
rect 18418 17176 18474 17232
rect 18326 15544 18382 15600
rect 18234 11192 18290 11248
rect 18602 18808 18658 18864
rect 18694 14864 18750 14920
rect 18510 12688 18566 12744
rect 18786 13096 18842 13152
rect 17958 7284 17960 7304
rect 17960 7284 18012 7304
rect 18012 7284 18014 7304
rect 17958 7248 18014 7284
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19246 19916 19302 19952
rect 19246 19896 19248 19916
rect 19248 19896 19300 19916
rect 19300 19896 19302 19916
rect 20626 21392 20682 21448
rect 19614 19760 19670 19816
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19522 18028 19524 18048
rect 19524 18028 19576 18048
rect 19576 18028 19578 18048
rect 19522 17992 19578 18028
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 18970 16088 19026 16144
rect 18878 12824 18934 12880
rect 18326 6296 18382 6352
rect 17958 4664 18014 4720
rect 18878 10104 18934 10160
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19062 15408 19118 15464
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19062 9560 19118 9616
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19614 13912 19670 13968
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19890 14456 19946 14512
rect 20350 18128 20406 18184
rect 20258 12144 20314 12200
rect 20902 16904 20958 16960
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 20626 16496 20682 16552
rect 20442 11600 20498 11656
rect 20442 9424 20498 9480
rect 20442 8880 20498 8936
rect 19890 6840 19946 6896
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21454 10648 21510 10704
rect 21178 9968 21234 10024
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21086 9152 21142 9208
rect 20994 8336 21050 8392
rect 21178 9016 21234 9072
rect 21362 8916 21364 8936
rect 21364 8916 21416 8936
rect 21416 8916 21418 8936
rect 21362 8880 21418 8916
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 21362 7928 21418 7984
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21270 7384 21326 7440
rect 21178 6704 21234 6760
rect 20442 5888 20498 5944
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21270 5072 21326 5128
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 18142 4120 18198 4176
rect 17958 4020 17960 4040
rect 17960 4020 18012 4040
rect 18012 4020 18014 4040
rect 17958 3984 18014 4020
rect 18050 3440 18106 3496
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17958 3052 18014 3088
rect 17958 3032 17960 3052
rect 17960 3032 18012 3052
rect 18012 3032 18014 3052
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 18970 2352 19026 2408
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19246 2524 19248 2544
rect 19248 2524 19300 2544
rect 19300 2524 19302 2544
rect 19246 2488 19302 2524
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 19154 1808 19210 1864
rect 19062 1400 19118 1456
<< metal3 >>
rect 20621 21450 20687 21453
rect 22200 21450 23000 21480
rect 20621 21448 23000 21450
rect 20621 21392 20626 21448
rect 20682 21392 23000 21448
rect 20621 21390 23000 21392
rect 20621 21387 20687 21390
rect 22200 21360 23000 21390
rect 17861 21042 17927 21045
rect 22200 21042 23000 21072
rect 17861 21040 23000 21042
rect 17861 20984 17866 21040
rect 17922 20984 23000 21040
rect 17861 20982 23000 20984
rect 17861 20979 17927 20982
rect 22200 20952 23000 20982
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 22200 20634 23000 20664
rect 22142 20544 23000 20634
rect 17953 20498 18019 20501
rect 22142 20498 22202 20544
rect 17953 20496 22202 20498
rect 17953 20440 17958 20496
rect 18014 20440 22202 20496
rect 17953 20438 22202 20440
rect 17953 20435 18019 20438
rect 22200 20226 23000 20256
rect 19566 20166 23000 20226
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 19241 19954 19307 19957
rect 19566 19954 19626 20166
rect 22200 20136 23000 20166
rect 19241 19952 19626 19954
rect 19241 19896 19246 19952
rect 19302 19896 19626 19952
rect 19241 19894 19626 19896
rect 19241 19891 19307 19894
rect 3877 19818 3943 19821
rect 19609 19818 19675 19821
rect 22200 19818 23000 19848
rect 3877 19816 19442 19818
rect 3877 19760 3882 19816
rect 3938 19760 19442 19816
rect 3877 19758 19442 19760
rect 3877 19755 3943 19758
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 19382 19410 19442 19758
rect 19609 19816 23000 19818
rect 19609 19760 19614 19816
rect 19670 19760 23000 19816
rect 19609 19758 23000 19760
rect 19609 19755 19675 19758
rect 22200 19728 23000 19758
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 22200 19410 23000 19440
rect 19382 19350 23000 19410
rect 22200 19320 23000 19350
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 22200 19002 23000 19032
rect 19566 18942 23000 19002
rect 18597 18866 18663 18869
rect 19566 18866 19626 18942
rect 22200 18912 23000 18942
rect 18597 18864 19626 18866
rect 18597 18808 18602 18864
rect 18658 18808 19626 18864
rect 18597 18806 19626 18808
rect 18597 18803 18663 18806
rect 18137 18730 18203 18733
rect 18137 18728 22202 18730
rect 18137 18672 18142 18728
rect 18198 18672 22202 18728
rect 18137 18670 22202 18672
rect 18137 18667 18203 18670
rect 22142 18624 22202 18670
rect 22142 18534 23000 18624
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 20345 18186 20411 18189
rect 22200 18186 23000 18216
rect 20345 18184 23000 18186
rect 20345 18128 20350 18184
rect 20406 18128 23000 18184
rect 20345 18126 23000 18128
rect 20345 18123 20411 18126
rect 22200 18096 23000 18126
rect 12341 18050 12407 18053
rect 13813 18050 13879 18053
rect 12341 18048 13879 18050
rect 12341 17992 12346 18048
rect 12402 17992 13818 18048
rect 13874 17992 13879 18048
rect 12341 17990 13879 17992
rect 12341 17987 12407 17990
rect 13813 17987 13879 17990
rect 19517 18052 19583 18053
rect 19517 18048 19564 18052
rect 19628 18050 19634 18052
rect 19517 17992 19522 18048
rect 19517 17988 19564 17992
rect 19628 17990 19674 18050
rect 19628 17988 19634 17990
rect 19517 17987 19583 17988
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 12249 17914 12315 17917
rect 13813 17914 13879 17917
rect 12249 17912 13879 17914
rect 12249 17856 12254 17912
rect 12310 17856 13818 17912
rect 13874 17856 13879 17912
rect 12249 17854 13879 17856
rect 12249 17851 12315 17854
rect 13813 17851 13879 17854
rect 17677 17778 17743 17781
rect 22200 17778 23000 17808
rect 17677 17776 23000 17778
rect 17677 17720 17682 17776
rect 17738 17720 23000 17776
rect 17677 17718 23000 17720
rect 17677 17715 17743 17718
rect 22200 17688 23000 17718
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 22200 17370 23000 17400
rect 22142 17280 23000 17370
rect 0 17234 800 17264
rect 3877 17234 3943 17237
rect 0 17232 3943 17234
rect 0 17176 3882 17232
rect 3938 17176 3943 17232
rect 0 17174 3943 17176
rect 0 17144 800 17174
rect 3877 17171 3943 17174
rect 18413 17234 18479 17237
rect 22142 17234 22202 17280
rect 18413 17232 22202 17234
rect 18413 17176 18418 17232
rect 18474 17176 22202 17232
rect 18413 17174 22202 17176
rect 18413 17171 18479 17174
rect 20897 16962 20963 16965
rect 22200 16962 23000 16992
rect 20897 16960 23000 16962
rect 20897 16904 20902 16960
rect 20958 16904 23000 16960
rect 20897 16902 23000 16904
rect 20897 16899 20963 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 20621 16554 20687 16557
rect 22200 16554 23000 16584
rect 20621 16552 23000 16554
rect 20621 16496 20626 16552
rect 20682 16496 23000 16552
rect 20621 16494 23000 16496
rect 20621 16491 20687 16494
rect 22200 16464 23000 16494
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 18965 16146 19031 16149
rect 22200 16146 23000 16176
rect 18965 16144 23000 16146
rect 18965 16088 18970 16144
rect 19026 16088 23000 16144
rect 18965 16086 23000 16088
rect 18965 16083 19031 16086
rect 22200 16056 23000 16086
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 22200 15738 23000 15768
rect 19566 15678 23000 15738
rect 18321 15602 18387 15605
rect 19566 15602 19626 15678
rect 22200 15648 23000 15678
rect 18321 15600 19626 15602
rect 18321 15544 18326 15600
rect 18382 15544 19626 15600
rect 18321 15542 19626 15544
rect 18321 15539 18387 15542
rect 19057 15466 19123 15469
rect 19057 15464 22202 15466
rect 19057 15408 19062 15464
rect 19118 15408 22202 15464
rect 19057 15406 22202 15408
rect 19057 15403 19123 15406
rect 22142 15360 22202 15406
rect 22142 15270 23000 15360
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 18689 14922 18755 14925
rect 22200 14922 23000 14952
rect 18689 14920 23000 14922
rect 18689 14864 18694 14920
rect 18750 14864 23000 14920
rect 18689 14862 23000 14864
rect 18689 14859 18755 14862
rect 22200 14832 23000 14862
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 19885 14514 19951 14517
rect 22200 14514 23000 14544
rect 19885 14512 23000 14514
rect 19885 14456 19890 14512
rect 19946 14456 23000 14512
rect 19885 14454 23000 14456
rect 19885 14451 19951 14454
rect 22200 14424 23000 14454
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 22200 14106 23000 14136
rect 22142 14016 23000 14106
rect 19609 13970 19675 13973
rect 22142 13970 22202 14016
rect 19609 13968 22202 13970
rect 19609 13912 19614 13968
rect 19670 13912 22202 13968
rect 19609 13910 22202 13912
rect 19609 13907 19675 13910
rect 22200 13698 23000 13728
rect 19566 13638 23000 13698
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 17953 13426 18019 13429
rect 19566 13426 19626 13638
rect 22200 13608 23000 13638
rect 17953 13424 19626 13426
rect 17953 13368 17958 13424
rect 18014 13368 19626 13424
rect 17953 13366 19626 13368
rect 17953 13363 18019 13366
rect 9581 13290 9647 13293
rect 19558 13290 19564 13292
rect 9581 13288 19564 13290
rect 9581 13232 9586 13288
rect 9642 13232 19564 13288
rect 9581 13230 19564 13232
rect 9581 13227 9647 13230
rect 19558 13228 19564 13230
rect 19628 13228 19634 13292
rect 22200 13290 23000 13320
rect 19750 13230 23000 13290
rect 18781 13154 18847 13157
rect 19750 13154 19810 13230
rect 22200 13200 23000 13230
rect 18781 13152 19810 13154
rect 18781 13096 18786 13152
rect 18842 13096 19810 13152
rect 18781 13094 19810 13096
rect 18781 13091 18847 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 18873 12882 18939 12885
rect 22200 12882 23000 12912
rect 18873 12880 23000 12882
rect 18873 12824 18878 12880
rect 18934 12824 23000 12880
rect 18873 12822 23000 12824
rect 18873 12819 18939 12822
rect 22200 12792 23000 12822
rect 18505 12746 18571 12749
rect 18505 12744 19626 12746
rect 18505 12688 18510 12744
rect 18566 12688 19626 12744
rect 18505 12686 19626 12688
rect 18505 12683 18571 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 19566 12474 19626 12686
rect 22200 12474 23000 12504
rect 19566 12414 23000 12474
rect 22200 12384 23000 12414
rect 20253 12202 20319 12205
rect 20253 12200 22202 12202
rect 20253 12144 20258 12200
rect 20314 12144 22202 12200
rect 20253 12142 22202 12144
rect 20253 12139 20319 12142
rect 22142 12096 22202 12142
rect 22142 12006 23000 12096
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 20437 11658 20503 11661
rect 22200 11658 23000 11688
rect 20437 11656 23000 11658
rect 20437 11600 20442 11656
rect 20498 11600 23000 11656
rect 20437 11598 23000 11600
rect 20437 11595 20503 11598
rect 22200 11568 23000 11598
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 12893 11250 12959 11253
rect 15285 11250 15351 11253
rect 12893 11248 15351 11250
rect 12893 11192 12898 11248
rect 12954 11192 15290 11248
rect 15346 11192 15351 11248
rect 12893 11190 15351 11192
rect 12893 11187 12959 11190
rect 15285 11187 15351 11190
rect 18229 11250 18295 11253
rect 22200 11250 23000 11280
rect 18229 11248 23000 11250
rect 18229 11192 18234 11248
rect 18290 11192 23000 11248
rect 18229 11190 23000 11192
rect 18229 11187 18295 11190
rect 22200 11160 23000 11190
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 22200 10842 23000 10872
rect 22142 10752 23000 10842
rect 21449 10706 21515 10709
rect 22142 10706 22202 10752
rect 21449 10704 22202 10706
rect 21449 10648 21454 10704
rect 21510 10648 22202 10704
rect 21449 10646 22202 10648
rect 21449 10643 21515 10646
rect 22200 10434 23000 10464
rect 19566 10374 23000 10434
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 18873 10162 18939 10165
rect 19566 10162 19626 10374
rect 22200 10344 23000 10374
rect 18873 10160 19626 10162
rect 18873 10104 18878 10160
rect 18934 10104 19626 10160
rect 18873 10102 19626 10104
rect 18873 10099 18939 10102
rect 21173 10026 21239 10029
rect 22200 10026 23000 10056
rect 21173 10024 23000 10026
rect 21173 9968 21178 10024
rect 21234 9968 23000 10024
rect 21173 9966 23000 9968
rect 21173 9963 21239 9966
rect 22200 9936 23000 9966
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 19057 9618 19123 9621
rect 22200 9618 23000 9648
rect 19057 9616 23000 9618
rect 19057 9560 19062 9616
rect 19118 9560 23000 9616
rect 19057 9558 23000 9560
rect 19057 9555 19123 9558
rect 22200 9528 23000 9558
rect 15837 9482 15903 9485
rect 20437 9482 20503 9485
rect 15837 9480 20503 9482
rect 15837 9424 15842 9480
rect 15898 9424 20442 9480
rect 20498 9424 20503 9480
rect 15837 9422 20503 9424
rect 15837 9419 15903 9422
rect 20437 9419 20503 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 21081 9210 21147 9213
rect 22200 9210 23000 9240
rect 21081 9208 23000 9210
rect 21081 9152 21086 9208
rect 21142 9152 23000 9208
rect 21081 9150 23000 9152
rect 21081 9147 21147 9150
rect 22200 9120 23000 9150
rect 15377 9074 15443 9077
rect 21173 9074 21239 9077
rect 15377 9072 21239 9074
rect 15377 9016 15382 9072
rect 15438 9016 21178 9072
rect 21234 9016 21239 9072
rect 15377 9014 21239 9016
rect 15377 9011 15443 9014
rect 21173 9011 21239 9014
rect 14181 8938 14247 8941
rect 15561 8938 15627 8941
rect 14181 8936 15627 8938
rect 14181 8880 14186 8936
rect 14242 8880 15566 8936
rect 15622 8880 15627 8936
rect 14181 8878 15627 8880
rect 14181 8875 14247 8878
rect 15561 8875 15627 8878
rect 15745 8938 15811 8941
rect 20437 8938 20503 8941
rect 15745 8936 20503 8938
rect 15745 8880 15750 8936
rect 15806 8880 20442 8936
rect 20498 8880 20503 8936
rect 15745 8878 20503 8880
rect 15745 8875 15811 8878
rect 20437 8875 20503 8878
rect 21357 8938 21423 8941
rect 21357 8936 22202 8938
rect 21357 8880 21362 8936
rect 21418 8880 22202 8936
rect 21357 8878 22202 8880
rect 21357 8875 21423 8878
rect 22142 8832 22202 8878
rect 22142 8742 23000 8832
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 20989 8394 21055 8397
rect 22200 8394 23000 8424
rect 20989 8392 23000 8394
rect 20989 8336 20994 8392
rect 21050 8336 23000 8392
rect 20989 8334 23000 8336
rect 20989 8331 21055 8334
rect 22200 8304 23000 8334
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 21357 7986 21423 7989
rect 22200 7986 23000 8016
rect 21357 7984 23000 7986
rect 21357 7928 21362 7984
rect 21418 7928 23000 7984
rect 21357 7926 23000 7928
rect 21357 7923 21423 7926
rect 22200 7896 23000 7926
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 22200 7578 23000 7608
rect 22142 7488 23000 7578
rect 21265 7442 21331 7445
rect 22142 7442 22202 7488
rect 21265 7440 22202 7442
rect 21265 7384 21270 7440
rect 21326 7384 22202 7440
rect 21265 7382 22202 7384
rect 21265 7379 21331 7382
rect 17953 7306 18019 7309
rect 17953 7304 19626 7306
rect 17953 7248 17958 7304
rect 18014 7248 19626 7304
rect 17953 7246 19626 7248
rect 17953 7243 18019 7246
rect 19566 7170 19626 7246
rect 22200 7170 23000 7200
rect 19566 7110 23000 7170
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 22200 7080 23000 7110
rect 19139 7039 19455 7040
rect 12617 6898 12683 6901
rect 19885 6898 19951 6901
rect 12617 6896 19951 6898
rect 12617 6840 12622 6896
rect 12678 6840 19890 6896
rect 19946 6840 19951 6896
rect 12617 6838 19951 6840
rect 12617 6835 12683 6838
rect 19885 6835 19951 6838
rect 21173 6762 21239 6765
rect 22200 6762 23000 6792
rect 21173 6760 23000 6762
rect 21173 6704 21178 6760
rect 21234 6704 23000 6760
rect 21173 6702 23000 6704
rect 21173 6699 21239 6702
rect 22200 6672 23000 6702
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 18321 6354 18387 6357
rect 22200 6354 23000 6384
rect 18321 6352 23000 6354
rect 18321 6296 18326 6352
rect 18382 6296 23000 6352
rect 18321 6294 23000 6296
rect 18321 6291 18387 6294
rect 22200 6264 23000 6294
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 20437 5946 20503 5949
rect 22200 5946 23000 5976
rect 20437 5944 23000 5946
rect 20437 5888 20442 5944
rect 20498 5888 23000 5944
rect 20437 5886 23000 5888
rect 20437 5883 20503 5886
rect 22200 5856 23000 5886
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 21590 5614 22202 5674
rect 17493 5538 17559 5541
rect 21590 5538 21650 5614
rect 17493 5536 21650 5538
rect 17493 5480 17498 5536
rect 17554 5480 21650 5536
rect 17493 5478 21650 5480
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 17493 5475 17559 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 6913 5266 6979 5269
rect 12709 5266 12775 5269
rect 6913 5264 12775 5266
rect 6913 5208 6918 5264
rect 6974 5208 12714 5264
rect 12770 5208 12775 5264
rect 6913 5206 12775 5208
rect 6913 5203 6979 5206
rect 12709 5203 12775 5206
rect 21265 5130 21331 5133
rect 22200 5130 23000 5160
rect 21265 5128 23000 5130
rect 21265 5072 21270 5128
rect 21326 5072 23000 5128
rect 21265 5070 23000 5072
rect 21265 5067 21331 5070
rect 22200 5040 23000 5070
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 17953 4722 18019 4725
rect 22200 4722 23000 4752
rect 17953 4720 23000 4722
rect 17953 4664 17958 4720
rect 18014 4664 23000 4720
rect 17953 4662 23000 4664
rect 17953 4659 18019 4662
rect 22200 4632 23000 4662
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 22200 4314 23000 4344
rect 22142 4224 23000 4314
rect 18137 4178 18203 4181
rect 22142 4178 22202 4224
rect 18137 4176 22202 4178
rect 18137 4120 18142 4176
rect 18198 4120 22202 4176
rect 18137 4118 22202 4120
rect 18137 4115 18203 4118
rect 17953 4042 18019 4045
rect 17953 4040 19626 4042
rect 17953 3984 17958 4040
rect 18014 3984 19626 4040
rect 17953 3982 19626 3984
rect 17953 3979 18019 3982
rect 19566 3906 19626 3982
rect 22200 3906 23000 3936
rect 19566 3846 23000 3906
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 18045 3498 18111 3501
rect 22200 3498 23000 3528
rect 18045 3496 23000 3498
rect 18045 3440 18050 3496
rect 18106 3440 23000 3496
rect 18045 3438 23000 3440
rect 18045 3435 18111 3438
rect 22200 3408 23000 3438
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 17953 3090 18019 3093
rect 22200 3090 23000 3120
rect 17953 3088 23000 3090
rect 17953 3032 17958 3088
rect 18014 3032 23000 3088
rect 17953 3030 23000 3032
rect 17953 3027 18019 3030
rect 22200 3000 23000 3030
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 22200 2682 23000 2712
rect 19566 2622 23000 2682
rect 19241 2546 19307 2549
rect 19566 2546 19626 2622
rect 22200 2592 23000 2622
rect 19241 2544 19626 2546
rect 19241 2488 19246 2544
rect 19302 2488 19626 2544
rect 19241 2486 19626 2488
rect 19241 2483 19307 2486
rect 18965 2410 19031 2413
rect 18965 2408 22202 2410
rect 18965 2352 18970 2408
rect 19026 2352 22202 2408
rect 18965 2350 22202 2352
rect 18965 2347 19031 2350
rect 22142 2304 22202 2350
rect 22142 2214 23000 2304
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 19149 1866 19215 1869
rect 22200 1866 23000 1896
rect 19149 1864 23000 1866
rect 19149 1808 19154 1864
rect 19210 1808 23000 1864
rect 19149 1806 23000 1808
rect 19149 1803 19215 1806
rect 22200 1776 23000 1806
rect 19057 1458 19123 1461
rect 22200 1458 23000 1488
rect 19057 1456 23000 1458
rect 19057 1400 19062 1456
rect 19118 1400 23000 1456
rect 19057 1398 23000 1400
rect 19057 1395 19123 1398
rect 22200 1368 23000 1398
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 19564 18048 19628 18052
rect 19564 17992 19578 18048
rect 19578 17992 19628 18048
rect 19564 17988 19628 17992
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 19564 13228 19628 13292
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 19563 18052 19629 18053
rect 19563 17988 19564 18052
rect 19628 17988 19629 18052
rect 19563 17987 19629 17988
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19566 13293 19626 17987
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 19563 13292 19629 13293
rect 19563 13228 19564 13292
rect 19628 13228 19629 13292
rect 19563 13227 19629 13228
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform -1 0 21344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform -1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform -1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform -1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform -1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform -1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1649977179
transform 1 0 19596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1649977179
transform -1 0 21344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1649977179
transform -1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1649977179
transform 1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 19596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 17296 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11960 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19688 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17112 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20608 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 17204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 12052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5796 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7268 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8096 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6164 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6348 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18400 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18676 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp 1649977179
transform 1 0 16008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1649977179
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_124
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_152
timestamp 1649977179
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1649977179
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_175
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_87
timestamp 1649977179
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1649977179
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_98
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_80
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_95
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1649977179
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_123
timestamp 1649977179
transform 1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_143
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_151
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_101
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_147
timestamp 1649977179
transform 1 0 14628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_171
timestamp 1649977179
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_183
timestamp 1649977179
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_84
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_97
timestamp 1649977179
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_126
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_154
timestamp 1649977179
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_211
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_119
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_131
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_160
timestamp 1649977179
transform 1 0 15824 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_172
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1649977179
transform 1 0 19596 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_207
timestamp 1649977179
transform 1 0 20148 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1649977179
transform 1 0 20516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1649977179
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_116
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_128
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_140
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_144
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1649977179
transform 1 0 18032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_213
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_218
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1649977179
transform 1 0 21528 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1649977179
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_96
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_106
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_118
timestamp 1649977179
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_199
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_216
timestamp 1649977179
transform 1 0 20976 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_220
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_78
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1649977179
transform 1 0 10672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1649977179
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1649977179
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_182
timestamp 1649977179
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_199
timestamp 1649977179
transform 1 0 19412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1649977179
transform 1 0 20148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_91
timestamp 1649977179
transform 1 0 9476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_103
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_152
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1649977179
transform 1 0 16100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1649977179
transform 1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_188
timestamp 1649977179
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1649977179
transform 1 0 19596 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1649977179
transform 1 0 20148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_213
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_85
timestamp 1649977179
transform 1 0 8924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_97
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_206
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_210
timestamp 1649977179
transform 1 0 20424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_68
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_95
timestamp 1649977179
transform 1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_104
timestamp 1649977179
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_68
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_79
timestamp 1649977179
transform 1 0 8372 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_83
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_92
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_133
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1649977179
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_187
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_191
timestamp 1649977179
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1649977179
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_181
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_213
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_66
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_78
timestamp 1649977179
transform 1 0 8280 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_90
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_102
timestamp 1649977179
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_192
timestamp 1649977179
transform 1 0 18768 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1649977179
transform 1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_214
timestamp 1649977179
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_218
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_54
timestamp 1649977179
transform 1 0 6072 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_66
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_100
timestamp 1649977179
transform 1 0 10304 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_112
timestamp 1649977179
transform 1 0 11408 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_124
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_135
timestamp 1649977179
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_49
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1649977179
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_69
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_94
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_98
timestamp 1649977179
transform 1 0 10120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_168
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_187
timestamp 1649977179
transform 1 0 18308 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1649977179
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_213
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_86
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1649977179
transform 1 0 9936 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_100
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_140
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_152
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_196
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1649977179
transform 1 0 20608 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_47
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_51
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_63
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1649977179
transform 1 0 7636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_92
timestamp 1649977179
transform 1 0 9568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1649977179
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1649977179
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_161
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1649977179
transform 1 0 17020 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_176
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_218
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_222
timestamp 1649977179
transform 1 0 21528 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1649977179
transform 1 0 7728 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_88
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_171
timestamp 1649977179
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_176
timestamp 1649977179
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_188
timestamp 1649977179
transform 1 0 18400 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1649977179
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_174
timestamp 1649977179
transform 1 0 17112 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_211
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1649977179
transform 1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_67
timestamp 1649977179
transform 1 0 7268 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_82
timestamp 1649977179
transform 1 0 8648 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_94
timestamp 1649977179
transform 1 0 9752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_183
timestamp 1649977179
transform 1 0 17940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_195
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1649977179
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_50
timestamp 1649977179
transform 1 0 5704 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1649977179
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_106
timestamp 1649977179
transform 1 0 10856 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_130
timestamp 1649977179
transform 1 0 13064 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1649977179
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 1649977179
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1649977179
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 1649977179
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_217
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_44
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1649977179
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_64
timestamp 1649977179
transform 1 0 6992 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_76
timestamp 1649977179
transform 1 0 8096 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_88
timestamp 1649977179
transform 1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_100
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_129
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_133
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_189
timestamp 1649977179
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1649977179
transform 1 0 20976 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1649977179
transform 1 0 6164 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_59
timestamp 1649977179
transform 1 0 6532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_95
timestamp 1649977179
transform 1 0 9844 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_99
timestamp 1649977179
transform 1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_103
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1649977179
transform 1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1649977179
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_176
timestamp 1649977179
transform 1 0 17296 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1649977179
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_41
timestamp 1649977179
transform 1 0 4876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1649977179
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_68
timestamp 1649977179
transform 1 0 7360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_73
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1649977179
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_100
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1649977179
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_138
timestamp 1649977179
transform 1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_154
timestamp 1649977179
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1649977179
transform 1 0 19504 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_204
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1649977179
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_35
timestamp 1649977179
transform 1 0 4324 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_45
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_57
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1649977179
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_91
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_95
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_143
timestamp 1649977179
transform 1 0 14260 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_149
timestamp 1649977179
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_170
timestamp 1649977179
transform 1 0 16744 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_199
timestamp 1649977179
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_203
timestamp 1649977179
transform 1 0 19780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_220
timestamp 1649977179
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_33
timestamp 1649977179
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1649977179
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1649977179
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_71
timestamp 1649977179
transform 1 0 7636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_91
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_98
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1649977179
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_129
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_133
timestamp 1649977179
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_145
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1649977179
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_196
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_200
timestamp 1649977179
transform 1 0 19504 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_216
timestamp 1649977179
transform 1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_45
timestamp 1649977179
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_70
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_91
timestamp 1649977179
transform 1 0 9476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_103
timestamp 1649977179
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_112
timestamp 1649977179
transform 1 0 11408 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_117
timestamp 1649977179
transform 1 0 11868 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1649977179
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1649977179
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_157
timestamp 1649977179
transform 1 0 15548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1649977179
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1649977179
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_201
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1649977179
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_91
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_96
timestamp 1649977179
transform 1 0 9936 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_176
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_188
timestamp 1649977179
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_206
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_210
timestamp 1649977179
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_216
timestamp 1649977179
transform 1 0 20976 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform 1 0 10028 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform 1 0 12144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1649977179
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1649977179
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1649977179
transform -1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1649977179
transform 1 0 7544 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1649977179
transform -1 0 5796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1649977179
transform -1 0 11776 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform 1 0 19688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform 1 0 14444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform 1 0 16928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform 1 0 4140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform -1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform -1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform -1 0 20148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform -1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform -1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform -1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform -1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform -1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1649977179
transform -1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1649977179
transform -1 0 21436 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1649977179
transform -1 0 21160 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1649977179
transform -1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1649977179
transform -1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1649977179
transform 1 0 17848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1649977179
transform -1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1649977179
transform -1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1649977179
transform -1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1649977179
transform -1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1649977179
transform -1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1649977179
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1649977179
transform -1 0 21160 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18768 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21252 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17388 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13156 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15088 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18308 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12788 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13064 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12144 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16284 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13340 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13340 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12144 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12328 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17756 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13064 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11592 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17296 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18032 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19872 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21252 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20976 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18768 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16928 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18308 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16652 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21344 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20424 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19320 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21252 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16100 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15088 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13892 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14812 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15824 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8280 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8372 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9660 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9476 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11224 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12236 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15180 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15272 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10580 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7360 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7728 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8280 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7360 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18216 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8280 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5244 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13064 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10488 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10028 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7636 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9752 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9476 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4968 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13340 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 16 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 17 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 18 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 19 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 20 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 21 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 22 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 23 nsew signal input
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 24 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 25 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 26 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 27 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 28 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 29 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 30 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 31 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 32 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 33 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 34 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 35 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 36 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 37 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 38 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 39 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 40 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 41 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 42 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 43 nsew signal tristate
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 44 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 45 nsew signal input
flabel metal2 s 7010 22200 7066 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 46 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 47 nsew signal input
flabel metal2 s 8114 22200 8170 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 48 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 49 nsew signal input
flabel metal2 s 9218 22200 9274 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 50 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 51 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 52 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 53 nsew signal input
flabel metal2 s 11426 22200 11482 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 54 nsew signal input
flabel metal2 s 1490 22200 1546 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 55 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 56 nsew signal input
flabel metal2 s 2594 22200 2650 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 57 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 58 nsew signal input
flabel metal2 s 3698 22200 3754 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 59 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 60 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 61 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 62 nsew signal input
flabel metal2 s 5906 22200 5962 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 63 nsew signal input
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 64 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 65 nsew signal tristate
flabel metal2 s 18050 22200 18106 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 66 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 67 nsew signal tristate
flabel metal2 s 19154 22200 19210 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 68 nsew signal tristate
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 69 nsew signal tristate
flabel metal2 s 20258 22200 20314 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 70 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 71 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 72 nsew signal tristate
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 73 nsew signal tristate
flabel metal2 s 22466 22200 22522 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 74 nsew signal tristate
flabel metal2 s 12530 22200 12586 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 75 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 76 nsew signal tristate
flabel metal2 s 13634 22200 13690 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 77 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 78 nsew signal tristate
flabel metal2 s 14738 22200 14794 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 79 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 80 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 81 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 82 nsew signal tristate
flabel metal2 s 16946 22200 17002 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 83 nsew signal tristate
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 84 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_11_
port 85 nsew signal input
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 right_bottom_grid_pin_13_
port 86 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 right_bottom_grid_pin_15_
port 87 nsew signal input
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 right_bottom_grid_pin_17_
port 88 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_1_
port 89 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_3_
port 90 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_5_
port 91 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_7_
port 92 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_9_
port 93 nsew signal input
flabel metal2 s 386 22200 442 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_1_
port 94 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
