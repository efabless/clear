magic
tech sky130A
magscale 1 2
timestamp 1656258101
<< viali >>
rect 3433 20553 3467 20587
rect 11989 20553 12023 20587
rect 12449 20553 12483 20587
rect 14289 20553 14323 20587
rect 15301 20553 15335 20587
rect 15853 20553 15887 20587
rect 16773 20553 16807 20587
rect 18429 20553 18463 20587
rect 19901 20553 19935 20587
rect 21097 20553 21131 20587
rect 1501 20485 1535 20519
rect 2145 20417 2179 20451
rect 2697 20417 2731 20451
rect 3249 20417 3283 20451
rect 3985 20417 4019 20451
rect 4445 20417 4479 20451
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 6009 20417 6043 20451
rect 6561 20417 6595 20451
rect 7021 20417 7055 20451
rect 7481 20417 7515 20451
rect 8125 20417 8159 20451
rect 8585 20417 8619 20451
rect 9321 20417 9355 20451
rect 10057 20417 10091 20451
rect 10701 20417 10735 20451
rect 10977 20417 11011 20451
rect 11805 20417 11839 20451
rect 12633 20417 12667 20451
rect 13277 20417 13311 20451
rect 14105 20417 14139 20451
rect 14657 20417 14691 20451
rect 15485 20417 15519 20451
rect 16037 20417 16071 20451
rect 16957 20417 16991 20451
rect 17509 20417 17543 20451
rect 18061 20417 18095 20451
rect 18613 20417 18647 20451
rect 19533 20417 19567 20451
rect 20085 20417 20119 20451
rect 20637 20417 20671 20451
rect 20913 20417 20947 20451
rect 1685 20349 1719 20383
rect 9045 20349 9079 20383
rect 9229 20349 9263 20383
rect 13001 20349 13035 20383
rect 13185 20349 13219 20383
rect 5549 20281 5583 20315
rect 7941 20281 7975 20315
rect 9689 20281 9723 20315
rect 10241 20281 10275 20315
rect 14841 20281 14875 20315
rect 17877 20281 17911 20315
rect 19349 20281 19383 20315
rect 20453 20281 20487 20315
rect 2329 20213 2363 20247
rect 2881 20213 2915 20247
rect 4169 20213 4203 20247
rect 4629 20213 4663 20247
rect 5089 20213 5123 20247
rect 5825 20213 5859 20247
rect 6745 20213 6779 20247
rect 7205 20213 7239 20247
rect 7665 20213 7699 20247
rect 8401 20213 8435 20247
rect 10517 20213 10551 20247
rect 11161 20213 11195 20247
rect 13645 20213 13679 20247
rect 17325 20213 17359 20247
rect 2053 20009 2087 20043
rect 2605 20009 2639 20043
rect 3065 20009 3099 20043
rect 3433 20009 3467 20043
rect 4537 20009 4571 20043
rect 5273 20009 5307 20043
rect 6285 20009 6319 20043
rect 9137 20009 9171 20043
rect 9413 20009 9447 20043
rect 13553 20009 13587 20043
rect 14197 20009 14231 20043
rect 14657 20009 14691 20043
rect 19441 20009 19475 20043
rect 4905 19941 4939 19975
rect 9873 19941 9907 19975
rect 15301 19941 15335 19975
rect 17141 19941 17175 19975
rect 5733 19873 5767 19907
rect 6653 19873 6687 19907
rect 6837 19873 6871 19907
rect 7757 19873 7791 19907
rect 12541 19873 12575 19907
rect 12909 19873 12943 19907
rect 13093 19873 13127 19907
rect 18429 19873 18463 19907
rect 18613 19873 18647 19907
rect 20269 19873 20303 19907
rect 1593 19805 1627 19839
rect 3801 19805 3835 19839
rect 8953 19805 8987 19839
rect 9597 19805 9631 19839
rect 10986 19805 11020 19839
rect 11253 19805 11287 19839
rect 11621 19805 11655 19839
rect 14381 19805 14415 19839
rect 14841 19805 14875 19839
rect 15117 19805 15151 19839
rect 15669 19805 15703 19839
rect 16129 19805 16163 19839
rect 16957 19805 16991 19839
rect 17693 19805 17727 19839
rect 18337 19805 18371 19839
rect 19257 19805 19291 19839
rect 21097 19805 21131 19839
rect 5825 19737 5859 19771
rect 16681 19737 16715 19771
rect 1777 19669 1811 19703
rect 3985 19669 4019 19703
rect 5917 19669 5951 19703
rect 6929 19669 6963 19703
rect 7297 19669 7331 19703
rect 7849 19669 7883 19703
rect 7941 19669 7975 19703
rect 8309 19669 8343 19703
rect 11805 19669 11839 19703
rect 13185 19669 13219 19703
rect 15853 19669 15887 19703
rect 16313 19669 16347 19703
rect 17509 19669 17543 19703
rect 17969 19669 18003 19703
rect 2237 19465 2271 19499
rect 4905 19465 4939 19499
rect 5273 19465 5307 19499
rect 6377 19465 6411 19499
rect 6929 19465 6963 19499
rect 7941 19465 7975 19499
rect 8585 19465 8619 19499
rect 9137 19465 9171 19499
rect 12909 19465 12943 19499
rect 17141 19465 17175 19499
rect 17601 19465 17635 19499
rect 18061 19465 18095 19499
rect 19625 19465 19659 19499
rect 20177 19465 20211 19499
rect 6009 19397 6043 19431
rect 7665 19397 7699 19431
rect 15178 19397 15212 19431
rect 1409 19329 1443 19363
rect 1869 19329 1903 19363
rect 4721 19329 4755 19363
rect 8401 19329 8435 19363
rect 9781 19329 9815 19363
rect 10037 19329 10071 19363
rect 14033 19329 14067 19363
rect 17417 19329 17451 19363
rect 17877 19329 17911 19363
rect 18337 19329 18371 19363
rect 18889 19329 18923 19363
rect 19441 19329 19475 19363
rect 19993 19329 20027 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 4261 19261 4295 19295
rect 14289 19261 14323 19295
rect 14933 19261 14967 19295
rect 9505 19193 9539 19227
rect 11161 19193 11195 19227
rect 18521 19193 18555 19227
rect 19073 19193 19107 19227
rect 1593 19125 1627 19159
rect 7297 19125 7331 19159
rect 11621 19125 11655 19159
rect 11897 19125 11931 19159
rect 12541 19125 12575 19159
rect 14565 19125 14599 19159
rect 16313 19125 16347 19159
rect 20729 19125 20763 19159
rect 21281 19125 21315 19159
rect 1409 18921 1443 18955
rect 7021 18921 7055 18955
rect 9045 18921 9079 18955
rect 10057 18921 10091 18955
rect 12449 18921 12483 18955
rect 18061 18921 18095 18955
rect 19349 18921 19383 18955
rect 6285 18853 6319 18887
rect 6653 18853 6687 18887
rect 17785 18853 17819 18887
rect 5641 18785 5675 18819
rect 5825 18785 5859 18819
rect 7481 18785 7515 18819
rect 7665 18785 7699 18819
rect 19809 18785 19843 18819
rect 5917 18717 5951 18751
rect 11713 18717 11747 18751
rect 17141 18717 17175 18751
rect 17601 18717 17635 18751
rect 18245 18717 18279 18751
rect 18613 18717 18647 18751
rect 19533 18717 19567 18751
rect 11446 18649 11480 18683
rect 20054 18649 20088 18683
rect 7389 18581 7423 18615
rect 8033 18581 8067 18615
rect 9689 18581 9723 18615
rect 10333 18581 10367 18615
rect 11989 18581 12023 18615
rect 13645 18581 13679 18615
rect 16497 18581 16531 18615
rect 16865 18581 16899 18615
rect 17325 18581 17359 18615
rect 18797 18581 18831 18615
rect 21189 18581 21223 18615
rect 7481 18377 7515 18411
rect 8493 18377 8527 18411
rect 19625 18377 19659 18411
rect 6745 18309 6779 18343
rect 10916 18309 10950 18343
rect 13062 18309 13096 18343
rect 17110 18309 17144 18343
rect 8401 18241 8435 18275
rect 12817 18241 12851 18275
rect 19165 18241 19199 18275
rect 19441 18241 19475 18275
rect 19993 18241 20027 18275
rect 20545 18241 20579 18275
rect 21097 18241 21131 18275
rect 5181 18173 5215 18207
rect 6469 18173 6503 18207
rect 6653 18173 6687 18207
rect 8677 18173 8711 18207
rect 11161 18173 11195 18207
rect 15945 18173 15979 18207
rect 16865 18173 16899 18207
rect 8033 18105 8067 18139
rect 9137 18105 9171 18139
rect 18613 18105 18647 18139
rect 20177 18105 20211 18139
rect 7113 18037 7147 18071
rect 9781 18037 9815 18071
rect 11621 18037 11655 18071
rect 14197 18037 14231 18071
rect 14473 18037 14507 18071
rect 18245 18037 18279 18071
rect 18981 18037 19015 18071
rect 20729 18037 20763 18071
rect 21281 18037 21315 18071
rect 4813 17833 4847 17867
rect 16221 17833 16255 17867
rect 17509 17833 17543 17867
rect 19717 17833 19751 17867
rect 5457 17697 5491 17731
rect 6653 17697 6687 17731
rect 7389 17697 7423 17731
rect 7481 17697 7515 17731
rect 8309 17697 8343 17731
rect 15669 17697 15703 17731
rect 18889 17697 18923 17731
rect 1685 17629 1719 17663
rect 5181 17629 5215 17663
rect 15853 17629 15887 17663
rect 16865 17629 16899 17663
rect 19257 17629 19291 17663
rect 21097 17629 21131 17663
rect 5273 17561 5307 17595
rect 7573 17561 7607 17595
rect 15761 17561 15795 17595
rect 18622 17561 18656 17595
rect 20830 17561 20864 17595
rect 1501 17493 1535 17527
rect 7941 17493 7975 17527
rect 17049 17493 17083 17527
rect 19441 17493 19475 17527
rect 5549 17289 5583 17323
rect 16037 17289 16071 17323
rect 16773 17289 16807 17323
rect 18797 17289 18831 17323
rect 19717 17289 19751 17323
rect 14136 17221 14170 17255
rect 10894 17153 10928 17187
rect 14913 17153 14947 17187
rect 19257 17153 19291 17187
rect 19533 17153 19567 17187
rect 19993 17153 20027 17187
rect 20545 17153 20579 17187
rect 21097 17153 21131 17187
rect 11161 17085 11195 17119
rect 14381 17085 14415 17119
rect 14657 17085 14691 17119
rect 19073 17017 19107 17051
rect 9781 16949 9815 16983
rect 11621 16949 11655 16983
rect 13001 16949 13035 16983
rect 20177 16949 20211 16983
rect 20729 16949 20763 16983
rect 21281 16949 21315 16983
rect 19625 16745 19659 16779
rect 18797 16677 18831 16711
rect 4813 16609 4847 16643
rect 6285 16609 6319 16643
rect 6929 16609 6963 16643
rect 7941 16609 7975 16643
rect 21005 16609 21039 16643
rect 21281 16609 21315 16643
rect 4905 16541 4939 16575
rect 4997 16541 5031 16575
rect 6101 16541 6135 16575
rect 10057 16541 10091 16575
rect 10313 16541 10347 16575
rect 11897 16541 11931 16575
rect 13553 16541 13587 16575
rect 14473 16541 14507 16575
rect 18153 16541 18187 16575
rect 18613 16541 18647 16575
rect 20749 16541 20783 16575
rect 8125 16473 8159 16507
rect 8953 16473 8987 16507
rect 12142 16473 12176 16507
rect 5365 16405 5399 16439
rect 5641 16405 5675 16439
rect 6009 16405 6043 16439
rect 7021 16405 7055 16439
rect 7113 16405 7147 16439
rect 7481 16405 7515 16439
rect 8033 16405 8067 16439
rect 8493 16405 8527 16439
rect 11437 16405 11471 16439
rect 13277 16405 13311 16439
rect 18337 16405 18371 16439
rect 5273 16201 5307 16235
rect 7297 16201 7331 16235
rect 8401 16201 8435 16235
rect 8861 16201 8895 16235
rect 15025 16201 15059 16235
rect 18981 16201 19015 16235
rect 19441 16201 19475 16235
rect 20269 16201 20303 16235
rect 13614 16133 13648 16167
rect 5365 16065 5399 16099
rect 8493 16065 8527 16099
rect 9137 16065 9171 16099
rect 17509 16065 17543 16099
rect 18153 16065 18187 16099
rect 18797 16065 18831 16099
rect 19257 16065 19291 16099
rect 19901 16065 19935 16099
rect 20545 16065 20579 16099
rect 21097 16065 21131 16099
rect 5181 15997 5215 16031
rect 8309 15997 8343 16031
rect 13369 15997 13403 16031
rect 5733 15929 5767 15963
rect 19717 15929 19751 15963
rect 6561 15861 6595 15895
rect 11529 15861 11563 15895
rect 14749 15861 14783 15895
rect 17693 15861 17727 15895
rect 18337 15861 18371 15895
rect 20729 15861 20763 15895
rect 21281 15861 21315 15895
rect 7665 15657 7699 15691
rect 12357 15657 12391 15691
rect 18429 15657 18463 15691
rect 19901 15657 19935 15691
rect 20545 15657 20579 15691
rect 5457 15521 5491 15555
rect 8125 15521 8159 15555
rect 8309 15521 8343 15555
rect 9781 15453 9815 15487
rect 11437 15453 11471 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 17049 15453 17083 15487
rect 18245 15453 18279 15487
rect 20085 15453 20119 15487
rect 20361 15453 20395 15487
rect 21097 15453 21131 15487
rect 10048 15385 10082 15419
rect 13470 15385 13504 15419
rect 16782 15385 16816 15419
rect 8033 15317 8067 15351
rect 8953 15317 8987 15351
rect 11161 15317 11195 15351
rect 15669 15317 15703 15351
rect 17417 15317 17451 15351
rect 21281 15317 21315 15351
rect 5549 15113 5583 15147
rect 6009 15113 6043 15147
rect 17141 15113 17175 15147
rect 20545 15113 20579 15147
rect 9934 15045 9968 15079
rect 5641 14977 5675 15011
rect 6377 14977 6411 15011
rect 9689 14977 9723 15011
rect 12642 14977 12676 15011
rect 16681 14977 16715 15011
rect 17325 14977 17359 15011
rect 20085 14977 20119 15011
rect 20729 14977 20763 15011
rect 21097 14977 21131 15011
rect 5457 14909 5491 14943
rect 7205 14909 7239 14943
rect 12909 14909 12943 14943
rect 11069 14841 11103 14875
rect 11529 14841 11563 14875
rect 16865 14841 16899 14875
rect 20269 14841 20303 14875
rect 13277 14773 13311 14807
rect 21281 14773 21315 14807
rect 7849 14569 7883 14603
rect 16865 14569 16899 14603
rect 19349 14569 19383 14603
rect 20269 14569 20303 14603
rect 7297 14433 7331 14467
rect 16037 14433 16071 14467
rect 16405 14433 16439 14467
rect 15770 14365 15804 14399
rect 16681 14365 16715 14399
rect 17325 14365 17359 14399
rect 20821 14365 20855 14399
rect 21097 14365 21131 14399
rect 7481 14297 7515 14331
rect 8125 14297 8159 14331
rect 17570 14297 17604 14331
rect 7389 14229 7423 14263
rect 11253 14229 11287 14263
rect 14657 14229 14691 14263
rect 18705 14229 18739 14263
rect 20637 14229 20671 14263
rect 21281 14229 21315 14263
rect 7113 14025 7147 14059
rect 7481 14025 7515 14059
rect 8309 14025 8343 14059
rect 9597 14025 9631 14059
rect 11529 14025 11563 14059
rect 12817 14025 12851 14059
rect 19257 14025 19291 14059
rect 20913 14025 20947 14059
rect 21189 14025 21223 14059
rect 10732 13957 10766 13991
rect 13952 13957 13986 13991
rect 18144 13957 18178 13991
rect 8125 13889 8159 13923
rect 10977 13889 11011 13923
rect 19533 13889 19567 13923
rect 19800 13889 19834 13923
rect 21373 13889 21407 13923
rect 6837 13821 6871 13855
rect 7021 13821 7055 13855
rect 14197 13821 14231 13855
rect 16773 13821 16807 13855
rect 17877 13821 17911 13855
rect 14565 13685 14599 13719
rect 7665 13481 7699 13515
rect 9965 13481 9999 13515
rect 11621 13481 11655 13515
rect 13461 13481 13495 13515
rect 16405 13481 16439 13515
rect 18889 13481 18923 13515
rect 19349 13481 19383 13515
rect 20637 13481 20671 13515
rect 21281 13481 21315 13515
rect 8125 13345 8159 13379
rect 8217 13345 8251 13379
rect 11345 13345 11379 13379
rect 12081 13345 12115 13379
rect 18061 13345 18095 13379
rect 14197 13277 14231 13311
rect 15025 13277 15059 13311
rect 15292 13277 15326 13311
rect 18521 13277 18555 13311
rect 19901 13277 19935 13311
rect 20361 13277 20395 13311
rect 20821 13277 20855 13311
rect 21097 13277 21131 13311
rect 8033 13209 8067 13243
rect 11078 13209 11112 13243
rect 12326 13209 12360 13243
rect 17794 13209 17828 13243
rect 9045 13141 9079 13175
rect 16681 13141 16715 13175
rect 18337 13141 18371 13175
rect 20177 13141 20211 13175
rect 7205 12937 7239 12971
rect 7665 12937 7699 12971
rect 11621 12937 11655 12971
rect 18521 12937 18555 12971
rect 20085 12937 20119 12971
rect 20729 12937 20763 12971
rect 21281 12937 21315 12971
rect 15761 12869 15795 12903
rect 7573 12801 7607 12835
rect 8677 12801 8711 12835
rect 10894 12801 10928 12835
rect 11161 12801 11195 12835
rect 14013 12801 14047 12835
rect 14280 12801 14314 12835
rect 16773 12801 16807 12835
rect 17040 12801 17074 12835
rect 20269 12801 20303 12835
rect 20545 12801 20579 12835
rect 21097 12801 21131 12835
rect 7849 12733 7883 12767
rect 8217 12733 8251 12767
rect 9781 12597 9815 12631
rect 15393 12597 15427 12631
rect 18153 12597 18187 12631
rect 19809 12597 19843 12631
rect 20269 12393 20303 12427
rect 20913 12393 20947 12427
rect 21189 12393 21223 12427
rect 19993 12325 20027 12359
rect 4905 12257 4939 12291
rect 6193 12257 6227 12291
rect 6377 12257 6411 12291
rect 7665 12257 7699 12291
rect 7849 12189 7883 12223
rect 10905 12189 10939 12223
rect 11161 12189 11195 12223
rect 15577 12189 15611 12223
rect 15853 12189 15887 12223
rect 19809 12189 19843 12223
rect 20453 12189 20487 12223
rect 20729 12189 20763 12223
rect 21373 12189 21407 12223
rect 4997 12121 5031 12155
rect 6101 12121 6135 12155
rect 6745 12121 6779 12155
rect 7757 12121 7791 12155
rect 15332 12121 15366 12155
rect 5089 12053 5123 12087
rect 5457 12053 5491 12087
rect 5733 12053 5767 12087
rect 8217 12053 8251 12087
rect 9781 12053 9815 12087
rect 11529 12053 11563 12087
rect 14197 12053 14231 12087
rect 19533 12053 19567 12087
rect 5549 11849 5583 11883
rect 7941 11849 7975 11883
rect 13921 11849 13955 11883
rect 21373 11849 21407 11883
rect 20760 11781 20794 11815
rect 7757 11713 7791 11747
rect 18521 11713 18555 11747
rect 21005 11645 21039 11679
rect 18797 11509 18831 11543
rect 19257 11509 19291 11543
rect 19625 11509 19659 11543
rect 11345 11305 11379 11339
rect 17325 11305 17359 11339
rect 21189 11305 21223 11339
rect 14105 11237 14139 11271
rect 20729 11237 20763 11271
rect 9965 11101 9999 11135
rect 11713 11101 11747 11135
rect 12357 11101 12391 11135
rect 15485 11101 15519 11135
rect 15761 11101 15795 11135
rect 18705 11101 18739 11135
rect 19349 11101 19383 11135
rect 21373 11101 21407 11135
rect 10232 11033 10266 11067
rect 12624 11033 12658 11067
rect 15218 11033 15252 11067
rect 18438 11033 18472 11067
rect 19594 11033 19628 11067
rect 13737 10965 13771 10999
rect 7389 10761 7423 10795
rect 19993 10761 20027 10795
rect 16948 10693 16982 10727
rect 7481 10625 7515 10659
rect 9689 10625 9723 10659
rect 9956 10625 9990 10659
rect 11621 10625 11655 10659
rect 11877 10625 11911 10659
rect 13369 10625 13403 10659
rect 13645 10625 13679 10659
rect 13901 10625 13935 10659
rect 19450 10625 19484 10659
rect 19717 10625 19751 10659
rect 21117 10625 21151 10659
rect 21373 10625 21407 10659
rect 7297 10557 7331 10591
rect 15393 10557 15427 10591
rect 16681 10557 16715 10591
rect 7849 10489 7883 10523
rect 18061 10489 18095 10523
rect 8125 10421 8159 10455
rect 11069 10421 11103 10455
rect 13001 10421 13035 10455
rect 15025 10421 15059 10455
rect 18337 10421 18371 10455
rect 11437 10217 11471 10251
rect 11805 10217 11839 10251
rect 16129 10217 16163 10251
rect 20085 10217 20119 10251
rect 11069 10149 11103 10183
rect 20821 10149 20855 10183
rect 9689 10081 9723 10115
rect 14749 10081 14783 10115
rect 18889 10013 18923 10047
rect 19901 10013 19935 10047
rect 20361 10013 20395 10047
rect 21005 10013 21039 10047
rect 9956 9945 9990 9979
rect 14994 9945 15028 9979
rect 16497 9945 16531 9979
rect 18245 9945 18279 9979
rect 19625 9945 19659 9979
rect 20545 9877 20579 9911
rect 21281 9877 21315 9911
rect 8217 9673 8251 9707
rect 19073 9673 19107 9707
rect 11529 9605 11563 9639
rect 18337 9605 18371 9639
rect 18705 9605 18739 9639
rect 8309 9537 8343 9571
rect 19349 9537 19383 9571
rect 19993 9537 20027 9571
rect 20269 9537 20303 9571
rect 20913 9537 20947 9571
rect 21189 9537 21223 9571
rect 8125 9469 8159 9503
rect 19533 9401 19567 9435
rect 20453 9401 20487 9435
rect 20729 9401 20763 9435
rect 21373 9401 21407 9435
rect 8677 9333 8711 9367
rect 15393 9333 15427 9367
rect 19809 9333 19843 9367
rect 8585 9129 8619 9163
rect 9413 9129 9447 9163
rect 11437 9129 11471 9163
rect 17693 9129 17727 9163
rect 19441 9129 19475 9163
rect 21097 9129 21131 9163
rect 13461 9061 13495 9095
rect 17417 9061 17451 9095
rect 8033 8993 8067 9027
rect 10517 8993 10551 9027
rect 10701 8993 10735 9027
rect 11989 8993 12023 9027
rect 12909 8993 12943 9027
rect 14565 8993 14599 9027
rect 14749 8993 14783 9027
rect 15669 8993 15703 9027
rect 15761 8993 15795 9027
rect 18337 8993 18371 9027
rect 19809 8993 19843 9027
rect 20637 8993 20671 9027
rect 17233 8925 17267 8959
rect 19257 8925 19291 8959
rect 20453 8925 20487 8959
rect 21281 8925 21315 8959
rect 8953 8857 8987 8891
rect 11897 8857 11931 8891
rect 15853 8857 15887 8891
rect 18061 8857 18095 8891
rect 18705 8857 18739 8891
rect 8125 8789 8159 8823
rect 8217 8789 8251 8823
rect 10793 8789 10827 8823
rect 11161 8789 11195 8823
rect 11805 8789 11839 8823
rect 13001 8789 13035 8823
rect 13093 8789 13127 8823
rect 14197 8789 14231 8823
rect 14841 8789 14875 8823
rect 15209 8789 15243 8823
rect 16221 8789 16255 8823
rect 18153 8789 18187 8823
rect 20085 8789 20119 8823
rect 20545 8789 20579 8823
rect 10425 8585 10459 8619
rect 12265 8585 12299 8619
rect 13185 8585 13219 8619
rect 13553 8585 13587 8619
rect 13645 8585 13679 8619
rect 14933 8585 14967 8619
rect 16221 8585 16255 8619
rect 16681 8585 16715 8619
rect 17141 8585 17175 8619
rect 18705 8585 18739 8619
rect 19533 8585 19567 8619
rect 20821 8585 20855 8619
rect 21281 8585 21315 8619
rect 11805 8517 11839 8551
rect 10793 8449 10827 8483
rect 11897 8449 11931 8483
rect 14197 8449 14231 8483
rect 16037 8449 16071 8483
rect 16865 8449 16899 8483
rect 17509 8449 17543 8483
rect 19441 8449 19475 8483
rect 20361 8449 20395 8483
rect 21005 8449 21039 8483
rect 10885 8381 10919 8415
rect 10977 8381 11011 8415
rect 11713 8381 11747 8415
rect 12633 8381 12667 8415
rect 13737 8381 13771 8415
rect 17601 8381 17635 8415
rect 17785 8381 17819 8415
rect 19625 8381 19659 8415
rect 14381 8313 14415 8347
rect 20545 8313 20579 8347
rect 19073 8245 19107 8279
rect 11713 8041 11747 8075
rect 17417 8041 17451 8075
rect 19625 8041 19659 8075
rect 20453 8041 20487 8075
rect 12081 7973 12115 8007
rect 14289 7973 14323 8007
rect 15577 7973 15611 8007
rect 20729 7973 20763 8007
rect 11253 7905 11287 7939
rect 17969 7905 18003 7939
rect 14105 7837 14139 7871
rect 15393 7837 15427 7871
rect 20269 7837 20303 7871
rect 20913 7837 20947 7871
rect 21373 7837 21407 7871
rect 17785 7769 17819 7803
rect 18429 7769 18463 7803
rect 19901 7769 19935 7803
rect 14657 7701 14691 7735
rect 17877 7701 17911 7735
rect 21189 7701 21223 7735
rect 19257 7497 19291 7531
rect 19993 7497 20027 7531
rect 21189 7497 21223 7531
rect 11989 7429 12023 7463
rect 18889 7429 18923 7463
rect 11069 7361 11103 7395
rect 19901 7361 19935 7395
rect 20545 7361 20579 7395
rect 21373 7361 21407 7395
rect 11805 7293 11839 7327
rect 11897 7293 11931 7327
rect 20085 7293 20119 7327
rect 19533 7225 19567 7259
rect 12357 7157 12391 7191
rect 15209 7157 15243 7191
rect 14657 6817 14691 6851
rect 15485 6817 15519 6851
rect 16589 6817 16623 6851
rect 17969 6817 18003 6851
rect 19809 6817 19843 6851
rect 21373 6817 21407 6851
rect 13461 6749 13495 6783
rect 16681 6749 16715 6783
rect 20361 6749 20395 6783
rect 21005 6749 21039 6783
rect 14565 6681 14599 6715
rect 16773 6681 16807 6715
rect 17877 6681 17911 6715
rect 18889 6681 18923 6715
rect 19625 6681 19659 6715
rect 13645 6613 13679 6647
rect 14105 6613 14139 6647
rect 14473 6613 14507 6647
rect 15669 6613 15703 6647
rect 15761 6613 15795 6647
rect 16129 6613 16163 6647
rect 17141 6613 17175 6647
rect 17417 6613 17451 6647
rect 17785 6613 17819 6647
rect 19257 6613 19291 6647
rect 19717 6613 19751 6647
rect 20545 6613 20579 6647
rect 20821 6613 20855 6647
rect 12265 6409 12299 6443
rect 13001 6409 13035 6443
rect 13461 6409 13495 6443
rect 14197 6409 14231 6443
rect 14933 6409 14967 6443
rect 15761 6409 15795 6443
rect 17417 6409 17451 6443
rect 17693 6409 17727 6443
rect 19533 6409 19567 6443
rect 20269 6409 20303 6443
rect 20637 6409 20671 6443
rect 21373 6409 21407 6443
rect 11069 6341 11103 6375
rect 11805 6341 11839 6375
rect 13093 6341 13127 6375
rect 17049 6341 17083 6375
rect 20729 6341 20763 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 11897 6273 11931 6307
rect 14105 6273 14139 6307
rect 18061 6273 18095 6307
rect 18889 6273 18923 6307
rect 19349 6273 19383 6307
rect 19809 6273 19843 6307
rect 11713 6205 11747 6239
rect 12909 6205 12943 6239
rect 14381 6205 14415 6239
rect 16865 6205 16899 6239
rect 16957 6205 16991 6239
rect 18153 6205 18187 6239
rect 18245 6205 18279 6239
rect 20821 6205 20855 6239
rect 1593 6137 1627 6171
rect 13737 6137 13771 6171
rect 16221 6137 16255 6171
rect 19073 6069 19107 6103
rect 19993 6069 20027 6103
rect 15117 5865 15151 5899
rect 17785 5865 17819 5899
rect 18797 5865 18831 5899
rect 19809 5865 19843 5899
rect 21281 5865 21315 5899
rect 20269 5797 20303 5831
rect 20729 5797 20763 5831
rect 15669 5729 15703 5763
rect 18337 5729 18371 5763
rect 19993 5661 20027 5695
rect 20453 5661 20487 5695
rect 20913 5661 20947 5695
rect 15485 5593 15519 5627
rect 16129 5593 16163 5627
rect 15577 5525 15611 5559
rect 18153 5525 18187 5559
rect 18245 5525 18279 5559
rect 19349 5525 19383 5559
rect 15117 5321 15151 5355
rect 19257 5321 19291 5355
rect 19625 5321 19659 5355
rect 21281 5321 21315 5355
rect 15485 5253 15519 5287
rect 19901 5185 19935 5219
rect 20545 5185 20579 5219
rect 20821 5185 20855 5219
rect 15577 5117 15611 5151
rect 15669 5117 15703 5151
rect 20361 5049 20395 5083
rect 21005 5049 21039 5083
rect 16129 4981 16163 5015
rect 18613 4981 18647 5015
rect 20085 4981 20119 5015
rect 19901 4777 19935 4811
rect 20637 4777 20671 4811
rect 20177 4709 20211 4743
rect 18153 4641 18187 4675
rect 19257 4573 19291 4607
rect 19717 4573 19751 4607
rect 20361 4573 20395 4607
rect 20821 4573 20855 4607
rect 17969 4505 18003 4539
rect 18613 4505 18647 4539
rect 21097 4505 21131 4539
rect 21281 4505 21315 4539
rect 17601 4437 17635 4471
rect 18061 4437 18095 4471
rect 19441 4437 19475 4471
rect 15209 4233 15243 4267
rect 17049 4233 17083 4267
rect 20269 4233 20303 4267
rect 20637 4233 20671 4267
rect 21281 4165 21315 4199
rect 15117 4097 15151 4131
rect 19901 4097 19935 4131
rect 14473 4029 14507 4063
rect 15025 4029 15059 4063
rect 16773 4029 16807 4063
rect 16957 4029 16991 4063
rect 21097 4029 21131 4063
rect 15577 3961 15611 3995
rect 17417 3961 17451 3995
rect 20177 3689 20211 3723
rect 20453 3689 20487 3723
rect 21097 3621 21131 3655
rect 19809 3417 19843 3451
rect 21281 3417 21315 3451
rect 21189 3145 21223 3179
rect 19349 3077 19383 3111
rect 20729 3077 20763 3111
rect 19717 3009 19751 3043
rect 20177 3009 20211 3043
rect 21281 3009 21315 3043
rect 18981 2941 19015 2975
rect 19993 2873 20027 2907
rect 20637 2805 20671 2839
rect 19993 2533 20027 2567
rect 20821 2465 20855 2499
rect 19349 2397 19383 2431
rect 20545 2397 20579 2431
rect 19717 2329 19751 2363
rect 20177 2329 20211 2363
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 3421 20587 3479 20593
rect 3421 20553 3433 20587
rect 3467 20584 3479 20587
rect 5626 20584 5632 20596
rect 3467 20556 5632 20584
rect 3467 20553 3479 20556
rect 3421 20547 3479 20553
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 10410 20584 10416 20596
rect 6932 20556 10416 20584
rect 382 20476 388 20528
rect 440 20516 446 20528
rect 1394 20516 1400 20528
rect 440 20488 1400 20516
rect 440 20476 446 20488
rect 1394 20476 1400 20488
rect 1452 20516 1458 20528
rect 1489 20519 1547 20525
rect 1489 20516 1501 20519
rect 1452 20488 1501 20516
rect 1452 20476 1458 20488
rect 1489 20485 1501 20488
rect 1535 20485 1547 20519
rect 5534 20516 5540 20528
rect 1489 20479 1547 20485
rect 5368 20488 5540 20516
rect 2038 20408 2044 20460
rect 2096 20448 2102 20460
rect 2133 20451 2191 20457
rect 2133 20448 2145 20451
rect 2096 20420 2145 20448
rect 2096 20408 2102 20420
rect 2133 20417 2145 20420
rect 2179 20417 2191 20451
rect 2133 20411 2191 20417
rect 2590 20408 2596 20460
rect 2648 20448 2654 20460
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2648 20420 2697 20448
rect 2648 20408 2654 20420
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 3142 20408 3148 20460
rect 3200 20448 3206 20460
rect 3237 20451 3295 20457
rect 3237 20448 3249 20451
rect 3200 20420 3249 20448
rect 3200 20408 3206 20420
rect 3237 20417 3249 20420
rect 3283 20417 3295 20451
rect 3237 20411 3295 20417
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20448 4031 20451
rect 4246 20448 4252 20460
rect 4019 20420 4252 20448
rect 4019 20417 4031 20420
rect 3973 20411 4031 20417
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4798 20448 4804 20460
rect 4479 20420 4804 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4798 20408 4804 20420
rect 4856 20408 4862 20460
rect 4893 20451 4951 20457
rect 4893 20417 4905 20451
rect 4939 20448 4951 20451
rect 5258 20448 5264 20460
rect 4939 20420 5264 20448
rect 4939 20417 4951 20420
rect 4893 20411 4951 20417
rect 5258 20408 5264 20420
rect 5316 20408 5322 20460
rect 5368 20457 5396 20488
rect 5534 20476 5540 20488
rect 5592 20516 5598 20528
rect 5902 20516 5908 20528
rect 5592 20488 5908 20516
rect 5592 20476 5598 20488
rect 5902 20476 5908 20488
rect 5960 20476 5966 20528
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20417 5411 20451
rect 5994 20448 6000 20460
rect 5907 20420 6000 20448
rect 5353 20411 5411 20417
rect 5994 20408 6000 20420
rect 6052 20448 6058 20460
rect 6454 20448 6460 20460
rect 6052 20420 6460 20448
rect 6052 20408 6058 20420
rect 6454 20408 6460 20420
rect 6512 20408 6518 20460
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 6638 20448 6644 20460
rect 6595 20420 6644 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 6638 20408 6644 20420
rect 6696 20448 6702 20460
rect 6822 20448 6828 20460
rect 6696 20420 6828 20448
rect 6696 20408 6702 20420
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20380 1731 20383
rect 6932 20380 6960 20556
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11974 20584 11980 20596
rect 11935 20556 11980 20584
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12526 20584 12532 20596
rect 12483 20556 12532 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 13136 20556 14289 20584
rect 13136 20544 13142 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15289 20587 15347 20593
rect 15289 20584 15301 20587
rect 14792 20556 15301 20584
rect 14792 20544 14798 20556
rect 15289 20553 15301 20556
rect 15335 20553 15347 20587
rect 15289 20547 15347 20553
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15436 20556 15853 20584
rect 15436 20544 15442 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 15930 20544 15936 20596
rect 15988 20584 15994 20596
rect 16761 20587 16819 20593
rect 16761 20584 16773 20587
rect 15988 20556 16773 20584
rect 15988 20544 15994 20556
rect 16761 20553 16773 20556
rect 16807 20553 16819 20587
rect 16761 20547 16819 20553
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 18417 20587 18475 20593
rect 18417 20584 18429 20587
rect 17552 20556 18429 20584
rect 17552 20544 17558 20556
rect 18417 20553 18429 20556
rect 18463 20553 18475 20587
rect 18417 20547 18475 20553
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19889 20587 19947 20593
rect 19889 20584 19901 20587
rect 19392 20556 19901 20584
rect 19392 20544 19398 20556
rect 19889 20553 19901 20556
rect 19935 20553 19947 20587
rect 19889 20547 19947 20553
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20312 20556 21097 20584
rect 20312 20544 20318 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 7558 20516 7564 20528
rect 7024 20488 7564 20516
rect 7024 20457 7052 20488
rect 7558 20476 7564 20488
rect 7616 20476 7622 20528
rect 9214 20476 9220 20528
rect 9272 20476 9278 20528
rect 19610 20516 19616 20528
rect 18616 20488 19616 20516
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7469 20451 7527 20457
rect 7469 20448 7481 20451
rect 7156 20420 7481 20448
rect 7156 20408 7162 20420
rect 7469 20417 7481 20420
rect 7515 20448 7527 20451
rect 8018 20448 8024 20460
rect 7515 20420 8024 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8202 20448 8208 20460
rect 8159 20420 8208 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 9232 20448 9260 20476
rect 8619 20420 9260 20448
rect 9309 20451 9367 20457
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9490 20448 9496 20460
rect 9355 20420 9496 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 9824 20420 10057 20448
rect 9824 20408 9830 20420
rect 10045 20417 10057 20420
rect 10091 20448 10103 20451
rect 10318 20448 10324 20460
rect 10091 20420 10324 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10686 20448 10692 20460
rect 10599 20420 10692 20448
rect 10686 20408 10692 20420
rect 10744 20448 10750 20460
rect 10870 20448 10876 20460
rect 10744 20420 10876 20448
rect 10744 20408 10750 20420
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20448 11023 20451
rect 11054 20448 11060 20460
rect 11011 20420 11060 20448
rect 11011 20417 11023 20420
rect 10965 20411 11023 20417
rect 11054 20408 11060 20420
rect 11112 20448 11118 20460
rect 11238 20448 11244 20460
rect 11112 20420 11244 20448
rect 11112 20408 11118 20420
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 1719 20352 6960 20380
rect 9033 20383 9091 20389
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 9033 20349 9045 20383
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 9398 20380 9404 20392
rect 9263 20352 9404 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 5537 20315 5595 20321
rect 5537 20281 5549 20315
rect 5583 20312 5595 20315
rect 6822 20312 6828 20324
rect 5583 20284 6828 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 6822 20272 6828 20284
rect 6880 20272 6886 20324
rect 7466 20272 7472 20324
rect 7524 20312 7530 20324
rect 7929 20315 7987 20321
rect 7929 20312 7941 20315
rect 7524 20284 7941 20312
rect 7524 20272 7530 20284
rect 7929 20281 7941 20284
rect 7975 20281 7987 20315
rect 7929 20275 7987 20281
rect 2314 20244 2320 20256
rect 2275 20216 2320 20244
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 2866 20244 2872 20256
rect 2827 20216 2872 20244
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 4154 20244 4160 20256
rect 4115 20216 4160 20244
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 4614 20244 4620 20256
rect 4575 20216 4620 20244
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 5077 20247 5135 20253
rect 5077 20213 5089 20247
rect 5123 20244 5135 20247
rect 5718 20244 5724 20256
rect 5123 20216 5724 20244
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 5810 20204 5816 20256
rect 5868 20244 5874 20256
rect 6730 20244 6736 20256
rect 5868 20216 5913 20244
rect 6691 20216 6736 20244
rect 5868 20204 5874 20216
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 7190 20244 7196 20256
rect 7151 20216 7196 20244
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 7650 20244 7656 20256
rect 7611 20216 7656 20244
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 8389 20247 8447 20253
rect 8389 20244 8401 20247
rect 7800 20216 8401 20244
rect 7800 20204 7806 20216
rect 8389 20213 8401 20216
rect 8435 20213 8447 20247
rect 9048 20244 9076 20343
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 11808 20380 11836 20411
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12584 20420 12633 20448
rect 12584 20408 12590 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12768 20420 13277 20448
rect 12768 20408 12774 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20417 14151 20451
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 14093 20411 14151 20417
rect 12986 20380 12992 20392
rect 9508 20352 11836 20380
rect 12947 20352 12992 20380
rect 9122 20272 9128 20324
rect 9180 20312 9186 20324
rect 9508 20312 9536 20352
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13538 20380 13544 20392
rect 13219 20352 13544 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13538 20340 13544 20352
rect 13596 20340 13602 20392
rect 9674 20312 9680 20324
rect 9180 20284 9536 20312
rect 9635 20284 9680 20312
rect 9180 20272 9186 20284
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 10229 20315 10287 20321
rect 10229 20281 10241 20315
rect 10275 20312 10287 20315
rect 13078 20312 13084 20324
rect 10275 20284 13084 20312
rect 10275 20281 10287 20284
rect 10229 20275 10287 20281
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 14108 20312 14136 20411
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15470 20448 15476 20460
rect 15431 20420 15476 20448
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20448 16083 20451
rect 16206 20448 16212 20460
rect 16071 20420 16212 20448
rect 16071 20417 16083 20420
rect 16025 20411 16083 20417
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20448 17003 20451
rect 17034 20448 17040 20460
rect 16991 20420 17040 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20448 17555 20451
rect 17586 20448 17592 20460
rect 17543 20420 17592 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 18046 20448 18052 20460
rect 18007 20420 18052 20448
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 18616 20457 18644 20488
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 21174 20516 21180 20528
rect 20088 20488 21180 20516
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20417 18659 20451
rect 18601 20411 18659 20417
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19886 20448 19892 20460
rect 19567 20420 19892 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 20088 20457 20116 20488
rect 21174 20476 21180 20488
rect 21232 20476 21238 20528
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20417 20683 20451
rect 20898 20448 20904 20460
rect 20859 20420 20904 20448
rect 20625 20411 20683 20417
rect 15286 20340 15292 20392
rect 15344 20380 15350 20392
rect 20640 20380 20668 20411
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 20990 20380 20996 20392
rect 15344 20352 19564 20380
rect 20640 20352 20996 20380
rect 15344 20340 15350 20352
rect 19536 20324 19564 20352
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 13188 20284 14136 20312
rect 9306 20244 9312 20256
rect 9048 20216 9312 20244
rect 8389 20207 8447 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 10502 20244 10508 20256
rect 10463 20216 10508 20244
rect 10502 20204 10508 20216
rect 10560 20204 10566 20256
rect 11149 20247 11207 20253
rect 11149 20213 11161 20247
rect 11195 20244 11207 20247
rect 12158 20244 12164 20256
rect 11195 20216 12164 20244
rect 11195 20213 11207 20216
rect 11149 20207 11207 20213
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 13188 20244 13216 20284
rect 14182 20272 14188 20324
rect 14240 20312 14246 20324
rect 14829 20315 14887 20321
rect 14829 20312 14841 20315
rect 14240 20284 14841 20312
rect 14240 20272 14246 20284
rect 14829 20281 14841 20284
rect 14875 20281 14887 20315
rect 14829 20275 14887 20281
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17865 20315 17923 20321
rect 17865 20312 17877 20315
rect 17000 20284 17877 20312
rect 17000 20272 17006 20284
rect 17865 20281 17877 20284
rect 17911 20281 17923 20315
rect 17865 20275 17923 20281
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 19337 20315 19395 20321
rect 19337 20312 19349 20315
rect 18196 20284 19349 20312
rect 18196 20272 18202 20284
rect 19337 20281 19349 20284
rect 19383 20281 19395 20315
rect 19337 20275 19395 20281
rect 19518 20272 19524 20324
rect 19576 20272 19582 20324
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 20441 20315 20499 20321
rect 20441 20312 20453 20315
rect 19760 20284 20453 20312
rect 19760 20272 19766 20284
rect 20441 20281 20453 20284
rect 20487 20281 20499 20315
rect 20441 20275 20499 20281
rect 12492 20216 13216 20244
rect 12492 20204 12498 20216
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13633 20247 13691 20253
rect 13633 20244 13645 20247
rect 13504 20216 13645 20244
rect 13504 20204 13510 20216
rect 13633 20213 13645 20216
rect 13679 20213 13691 20247
rect 13633 20207 13691 20213
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17313 20247 17371 20253
rect 17313 20244 17325 20247
rect 16632 20216 17325 20244
rect 16632 20204 16638 20216
rect 17313 20213 17325 20216
rect 17359 20213 17371 20247
rect 17313 20207 17371 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 2590 20040 2596 20052
rect 2551 20012 2596 20040
rect 2590 20000 2596 20012
rect 2648 20000 2654 20052
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20040 3111 20043
rect 3142 20040 3148 20052
rect 3099 20012 3148 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 3142 20000 3148 20012
rect 3200 20000 3206 20052
rect 3418 20040 3424 20052
rect 3379 20012 3424 20040
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 4798 20040 4804 20052
rect 4571 20012 4804 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20040 5319 20043
rect 5994 20040 6000 20052
rect 5307 20012 6000 20040
rect 5307 20009 5319 20012
rect 5261 20003 5319 20009
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6273 20043 6331 20049
rect 6273 20009 6285 20043
rect 6319 20040 6331 20043
rect 9122 20040 9128 20052
rect 6319 20012 8984 20040
rect 9083 20012 9128 20040
rect 6319 20009 6331 20012
rect 6273 20003 6331 20009
rect 4893 19975 4951 19981
rect 4893 19941 4905 19975
rect 4939 19972 4951 19975
rect 5534 19972 5540 19984
rect 4939 19944 5540 19972
rect 4939 19941 4951 19944
rect 4893 19935 4951 19941
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 8846 19972 8852 19984
rect 5736 19944 8852 19972
rect 5736 19913 5764 19944
rect 8846 19932 8852 19944
rect 8904 19932 8910 19984
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19873 6699 19907
rect 6822 19904 6828 19916
rect 6783 19876 6828 19904
rect 6641 19867 6699 19873
rect 1486 19796 1492 19848
rect 1544 19836 1550 19848
rect 1581 19839 1639 19845
rect 1581 19836 1593 19839
rect 1544 19808 1593 19836
rect 1544 19796 1550 19808
rect 1581 19805 1593 19808
rect 1627 19805 1639 19839
rect 1581 19799 1639 19805
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 3476 19808 3801 19836
rect 3476 19796 3482 19808
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 6656 19836 6684 19867
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7745 19907 7803 19913
rect 6932 19876 7696 19904
rect 6932 19836 6960 19876
rect 6656 19808 6960 19836
rect 7668 19836 7696 19876
rect 7745 19873 7757 19907
rect 7791 19904 7803 19907
rect 8018 19904 8024 19916
rect 7791 19876 8024 19904
rect 7791 19873 7803 19876
rect 7745 19867 7803 19873
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8956 19904 8984 20012
rect 9122 20000 9128 20012
rect 9180 20000 9186 20052
rect 9398 20040 9404 20052
rect 9359 20012 9404 20040
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 13538 20040 13544 20052
rect 9508 20012 12434 20040
rect 13499 20012 13544 20040
rect 9030 19932 9036 19984
rect 9088 19972 9094 19984
rect 9508 19972 9536 20012
rect 9858 19972 9864 19984
rect 9088 19944 9536 19972
rect 9819 19944 9864 19972
rect 9088 19932 9094 19944
rect 9858 19932 9864 19944
rect 9916 19932 9922 19984
rect 8956 19876 9720 19904
rect 7668 19808 8616 19836
rect 3789 19799 3847 19805
rect 5813 19771 5871 19777
rect 5813 19737 5825 19771
rect 5859 19768 5871 19771
rect 7006 19768 7012 19780
rect 5859 19740 7012 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 7374 19768 7380 19780
rect 7208 19740 7380 19768
rect 1762 19700 1768 19712
rect 1723 19672 1768 19700
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 3970 19700 3976 19712
rect 3931 19672 3976 19700
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 5902 19660 5908 19712
rect 5960 19700 5966 19712
rect 6917 19703 6975 19709
rect 5960 19672 6005 19700
rect 5960 19660 5966 19672
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7208 19700 7236 19740
rect 7374 19728 7380 19740
rect 7432 19728 7438 19780
rect 6963 19672 7236 19700
rect 7285 19703 7343 19709
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7285 19669 7297 19703
rect 7331 19700 7343 19703
rect 7837 19703 7895 19709
rect 7837 19700 7849 19703
rect 7331 19672 7849 19700
rect 7331 19669 7343 19672
rect 7285 19663 7343 19669
rect 7837 19669 7849 19672
rect 7883 19669 7895 19703
rect 7837 19663 7895 19669
rect 7926 19660 7932 19712
rect 7984 19700 7990 19712
rect 8297 19703 8355 19709
rect 7984 19672 8029 19700
rect 7984 19660 7990 19672
rect 8297 19669 8309 19703
rect 8343 19700 8355 19703
rect 8478 19700 8484 19712
rect 8343 19672 8484 19700
rect 8343 19669 8355 19672
rect 8297 19663 8355 19669
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 8588 19700 8616 19808
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8720 19808 8953 19836
rect 8720 19796 8726 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 9582 19836 9588 19848
rect 9543 19808 9588 19836
rect 8941 19799 8999 19805
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 9692 19768 9720 19876
rect 10962 19796 10968 19848
rect 11020 19845 11026 19848
rect 11020 19836 11032 19845
rect 11238 19836 11244 19848
rect 11020 19808 11065 19836
rect 11199 19808 11244 19836
rect 11020 19799 11032 19808
rect 11020 19796 11026 19799
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11609 19839 11667 19845
rect 11609 19805 11621 19839
rect 11655 19805 11667 19839
rect 12406 19836 12434 20012
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 13872 20012 14197 20040
rect 13872 20000 13878 20012
rect 14185 20009 14197 20012
rect 14231 20009 14243 20043
rect 14642 20040 14648 20052
rect 14603 20012 14648 20040
rect 14185 20003 14243 20009
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 17862 20040 17868 20052
rect 14752 20012 17868 20040
rect 14752 19972 14780 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18598 20000 18604 20052
rect 18656 20040 18662 20052
rect 19429 20043 19487 20049
rect 19429 20040 19441 20043
rect 18656 20012 19441 20040
rect 18656 20000 18662 20012
rect 19429 20009 19441 20012
rect 19475 20009 19487 20043
rect 19429 20003 19487 20009
rect 15286 19972 15292 19984
rect 12820 19944 14780 19972
rect 15247 19944 15292 19972
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19904 12587 19907
rect 12710 19904 12716 19916
rect 12575 19876 12716 19904
rect 12575 19873 12587 19876
rect 12529 19867 12587 19873
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 12618 19836 12624 19848
rect 12406 19808 12624 19836
rect 11609 19799 11667 19805
rect 11624 19768 11652 19799
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 9692 19740 11652 19768
rect 11698 19728 11704 19780
rect 11756 19768 11762 19780
rect 12434 19768 12440 19780
rect 11756 19740 12440 19768
rect 11756 19728 11762 19740
rect 12434 19728 12440 19740
rect 12492 19728 12498 19780
rect 11146 19700 11152 19712
rect 8588 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11793 19703 11851 19709
rect 11793 19669 11805 19703
rect 11839 19700 11851 19703
rect 12820 19700 12848 19944
rect 15286 19932 15292 19944
rect 15344 19932 15350 19984
rect 17129 19975 17187 19981
rect 17129 19941 17141 19975
rect 17175 19972 17187 19975
rect 17175 19944 19288 19972
rect 17175 19941 17187 19944
rect 17129 19935 17187 19941
rect 12897 19907 12955 19913
rect 12897 19873 12909 19907
rect 12943 19873 12955 19907
rect 13078 19904 13084 19916
rect 13039 19876 13084 19904
rect 12897 19867 12955 19873
rect 12912 19836 12940 19867
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 13446 19864 13452 19916
rect 13504 19904 13510 19916
rect 13504 19876 15700 19904
rect 13504 19864 13510 19876
rect 14369 19839 14427 19845
rect 12912 19808 14320 19836
rect 14292 19768 14320 19808
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14458 19836 14464 19848
rect 14415 19808 14464 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14826 19836 14832 19848
rect 14787 19808 14832 19836
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 15102 19836 15108 19848
rect 15063 19808 15108 19836
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 15672 19845 15700 19876
rect 17218 19864 17224 19916
rect 17276 19904 17282 19916
rect 17276 19876 18368 19904
rect 17276 19864 17282 19876
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 16114 19836 16120 19848
rect 16075 19808 16120 19836
rect 15657 19799 15715 19805
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 17126 19836 17132 19848
rect 16991 19808 17132 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 18340 19845 18368 19876
rect 18414 19864 18420 19916
rect 18472 19904 18478 19916
rect 18598 19904 18604 19916
rect 18472 19876 18517 19904
rect 18559 19876 18604 19904
rect 18472 19864 18478 19876
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 19260 19845 19288 19944
rect 19794 19864 19800 19916
rect 19852 19904 19858 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 19852 19876 20269 19904
rect 19852 19864 19858 19876
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 20257 19867 20315 19873
rect 18325 19839 18383 19845
rect 18325 19805 18337 19839
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 21082 19836 21088 19848
rect 21043 19808 21088 19836
rect 19245 19799 19303 19805
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 16390 19768 16396 19780
rect 14292 19740 16396 19768
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 16669 19771 16727 19777
rect 16669 19737 16681 19771
rect 16715 19768 16727 19771
rect 21100 19768 21128 19796
rect 16715 19740 21128 19768
rect 16715 19737 16727 19740
rect 16669 19731 16727 19737
rect 13170 19700 13176 19712
rect 11839 19672 12848 19700
rect 13131 19672 13176 19700
rect 11839 19669 11851 19672
rect 11793 19663 11851 19669
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 15838 19700 15844 19712
rect 15799 19672 15844 19700
rect 15838 19660 15844 19672
rect 15896 19660 15902 19712
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 17402 19700 17408 19712
rect 16347 19672 17408 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 17770 19700 17776 19712
rect 17543 19672 17776 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 17770 19660 17776 19672
rect 17828 19660 17834 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18230 19700 18236 19712
rect 18003 19672 18236 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 2225 19499 2283 19505
rect 2225 19496 2237 19499
rect 1544 19468 2237 19496
rect 1544 19456 1550 19468
rect 2225 19465 2237 19468
rect 2271 19465 2283 19499
rect 2225 19459 2283 19465
rect 4893 19499 4951 19505
rect 4893 19465 4905 19499
rect 4939 19465 4951 19499
rect 5258 19496 5264 19508
rect 5219 19468 5264 19496
rect 4893 19459 4951 19465
rect 4908 19428 4936 19459
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 5902 19456 5908 19508
rect 5960 19496 5966 19508
rect 6365 19499 6423 19505
rect 6365 19496 6377 19499
rect 5960 19468 6377 19496
rect 5960 19456 5966 19468
rect 6365 19465 6377 19468
rect 6411 19465 6423 19499
rect 6365 19459 6423 19465
rect 6917 19499 6975 19505
rect 6917 19465 6929 19499
rect 6963 19496 6975 19499
rect 7098 19496 7104 19508
rect 6963 19468 7104 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 7926 19496 7932 19508
rect 7887 19468 7932 19496
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8573 19499 8631 19505
rect 8076 19468 8524 19496
rect 8076 19456 8082 19468
rect 5997 19431 6055 19437
rect 4908 19400 5948 19428
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19360 1455 19363
rect 1857 19363 1915 19369
rect 1857 19360 1869 19363
rect 1443 19332 1869 19360
rect 1443 19329 1455 19332
rect 1397 19323 1455 19329
rect 1857 19329 1869 19332
rect 1903 19329 1915 19363
rect 4706 19360 4712 19372
rect 4667 19332 4712 19360
rect 1857 19323 1915 19329
rect 934 19252 940 19304
rect 992 19292 998 19304
rect 1412 19292 1440 19323
rect 4706 19320 4712 19332
rect 4764 19320 4770 19372
rect 5920 19360 5948 19400
rect 5997 19397 6009 19431
rect 6043 19428 6055 19431
rect 6638 19428 6644 19440
rect 6043 19400 6644 19428
rect 6043 19397 6055 19400
rect 5997 19391 6055 19397
rect 6638 19388 6644 19400
rect 6696 19388 6702 19440
rect 7653 19431 7711 19437
rect 7653 19397 7665 19431
rect 7699 19428 7711 19431
rect 8202 19428 8208 19440
rect 7699 19400 8208 19428
rect 7699 19397 7711 19400
rect 7653 19391 7711 19397
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 6914 19360 6920 19372
rect 5920 19332 6920 19360
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 8389 19363 8447 19369
rect 8389 19360 8401 19363
rect 8352 19332 8401 19360
rect 8352 19320 8358 19332
rect 8389 19329 8401 19332
rect 8435 19329 8447 19363
rect 8496 19360 8524 19468
rect 8573 19465 8585 19499
rect 8619 19465 8631 19499
rect 8573 19459 8631 19465
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 9582 19496 9588 19508
rect 9171 19468 9588 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 8588 19428 8616 19459
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 11698 19496 11704 19508
rect 9692 19468 11704 19496
rect 9692 19428 9720 19468
rect 11698 19456 11704 19468
rect 11756 19456 11762 19508
rect 11790 19456 11796 19508
rect 11848 19496 11854 19508
rect 12897 19499 12955 19505
rect 12897 19496 12909 19499
rect 11848 19468 12909 19496
rect 11848 19456 11854 19468
rect 12897 19465 12909 19468
rect 12943 19465 12955 19499
rect 12897 19459 12955 19465
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17218 19496 17224 19508
rect 17175 19468 17224 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17589 19499 17647 19505
rect 17589 19465 17601 19499
rect 17635 19465 17647 19499
rect 17589 19459 17647 19465
rect 18049 19499 18107 19505
rect 18049 19465 18061 19499
rect 18095 19496 18107 19499
rect 19610 19496 19616 19508
rect 18095 19468 19472 19496
rect 19571 19468 19616 19496
rect 18095 19465 18107 19468
rect 18049 19459 18107 19465
rect 11238 19428 11244 19440
rect 8588 19400 9720 19428
rect 9784 19400 11244 19428
rect 9674 19360 9680 19372
rect 8496 19332 9680 19360
rect 8389 19323 8447 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 9784 19369 9812 19400
rect 11238 19388 11244 19400
rect 11296 19428 11302 19440
rect 11882 19428 11888 19440
rect 11296 19400 11888 19428
rect 11296 19388 11302 19400
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 15166 19431 15224 19437
rect 15166 19428 15178 19431
rect 12676 19400 15178 19428
rect 12676 19388 12682 19400
rect 15166 19397 15178 19400
rect 15212 19428 15224 19431
rect 16022 19428 16028 19440
rect 15212 19400 16028 19428
rect 15212 19397 15224 19400
rect 15166 19391 15224 19397
rect 16022 19388 16028 19400
rect 16080 19388 16086 19440
rect 17604 19428 17632 19459
rect 17604 19400 18368 19428
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19329 9827 19363
rect 9769 19323 9827 19329
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 10025 19363 10083 19369
rect 10025 19360 10037 19363
rect 9916 19332 10037 19360
rect 9916 19320 9922 19332
rect 10025 19329 10037 19332
rect 10071 19329 10083 19363
rect 10025 19323 10083 19329
rect 11146 19320 11152 19372
rect 11204 19360 11210 19372
rect 12710 19360 12716 19372
rect 11204 19332 12716 19360
rect 11204 19320 11210 19332
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 14021 19363 14079 19369
rect 14021 19360 14033 19363
rect 13044 19332 14033 19360
rect 13044 19320 13050 19332
rect 14021 19329 14033 19332
rect 14067 19360 14079 19363
rect 17405 19363 17463 19369
rect 14067 19332 17356 19360
rect 14067 19329 14079 19332
rect 14021 19323 14079 19329
rect 4246 19292 4252 19304
rect 992 19264 1440 19292
rect 4207 19264 4252 19292
rect 992 19252 998 19264
rect 4246 19252 4252 19264
rect 4304 19252 4310 19304
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 9876 19292 9904 19320
rect 8260 19264 9904 19292
rect 8260 19252 8266 19264
rect 9493 19227 9551 19233
rect 9493 19193 9505 19227
rect 9539 19224 9551 19227
rect 9766 19224 9772 19236
rect 9539 19196 9772 19224
rect 9539 19193 9551 19196
rect 9493 19187 9551 19193
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 11164 19233 11192 19320
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14323 19264 14933 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 11149 19227 11207 19233
rect 11149 19193 11161 19227
rect 11195 19193 11207 19227
rect 12066 19224 12072 19236
rect 11149 19187 11207 19193
rect 11256 19196 12072 19224
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 7285 19159 7343 19165
rect 7285 19125 7297 19159
rect 7331 19156 7343 19159
rect 7374 19156 7380 19168
rect 7331 19128 7380 19156
rect 7331 19125 7343 19128
rect 7285 19119 7343 19125
rect 7374 19116 7380 19128
rect 7432 19156 7438 19168
rect 11256 19156 11284 19196
rect 12066 19184 12072 19196
rect 12124 19184 12130 19236
rect 14384 19168 14412 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 17328 19224 17356 19332
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 17451 19332 17816 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 17788 19292 17816 19332
rect 17862 19320 17868 19372
rect 17920 19360 17926 19372
rect 18340 19369 18368 19400
rect 18325 19363 18383 19369
rect 17920 19332 17965 19360
rect 17920 19320 17926 19332
rect 18325 19329 18337 19363
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 18506 19320 18512 19372
rect 18564 19320 18570 19372
rect 18874 19360 18880 19372
rect 18835 19332 18880 19360
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19058 19320 19064 19372
rect 19116 19320 19122 19372
rect 19444 19369 19472 19468
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19496 20223 19499
rect 20622 19496 20628 19508
rect 20211 19468 20628 19496
rect 20211 19465 20223 19468
rect 20165 19459 20223 19465
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 19536 19400 20576 19428
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 18046 19292 18052 19304
rect 17788 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 17954 19224 17960 19236
rect 17328 19196 17960 19224
rect 17954 19184 17960 19196
rect 18012 19184 18018 19236
rect 18524 19233 18552 19320
rect 19076 19233 19104 19320
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19536 19292 19564 19400
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20548 19369 20576 19400
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 20806 19320 20812 19372
rect 20864 19360 20870 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20864 19332 21097 19360
rect 20864 19320 20870 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 19208 19264 19564 19292
rect 19208 19252 19214 19264
rect 18509 19227 18567 19233
rect 18509 19193 18521 19227
rect 18555 19193 18567 19227
rect 18509 19187 18567 19193
rect 19061 19227 19119 19233
rect 19061 19193 19073 19227
rect 19107 19193 19119 19227
rect 19061 19187 19119 19193
rect 7432 19128 11284 19156
rect 11609 19159 11667 19165
rect 7432 19116 7438 19128
rect 11609 19125 11621 19159
rect 11655 19156 11667 19159
rect 11882 19156 11888 19168
rect 11655 19128 11888 19156
rect 11655 19125 11667 19128
rect 11609 19119 11667 19125
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12526 19156 12532 19168
rect 12487 19128 12532 19156
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 14366 19116 14372 19168
rect 14424 19156 14430 19168
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 14424 19128 14565 19156
rect 14424 19116 14430 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 14553 19119 14611 19125
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19156 16359 19159
rect 17218 19156 17224 19168
rect 16347 19128 17224 19156
rect 16347 19125 16359 19128
rect 16301 19119 16359 19125
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1394 18952 1400 18964
rect 1355 18924 1400 18952
rect 1394 18912 1400 18924
rect 1452 18912 1458 18964
rect 7006 18952 7012 18964
rect 6967 18924 7012 18952
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 9033 18955 9091 18961
rect 9033 18921 9045 18955
rect 9079 18952 9091 18955
rect 9214 18952 9220 18964
rect 9079 18924 9220 18952
rect 9079 18921 9091 18924
rect 9033 18915 9091 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10686 18952 10692 18964
rect 10091 18924 10692 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 11112 18924 12449 18952
rect 11112 18912 11118 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 18046 18952 18052 18964
rect 18007 18924 18052 18952
rect 12437 18915 12495 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19337 18955 19395 18961
rect 19337 18921 19349 18955
rect 19383 18952 19395 18955
rect 21358 18952 21364 18964
rect 19383 18924 21364 18952
rect 19383 18921 19395 18924
rect 19337 18915 19395 18921
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 6273 18887 6331 18893
rect 6273 18853 6285 18887
rect 6319 18884 6331 18887
rect 6546 18884 6552 18896
rect 6319 18856 6552 18884
rect 6319 18853 6331 18856
rect 6273 18847 6331 18853
rect 6546 18844 6552 18856
rect 6604 18844 6610 18896
rect 6641 18887 6699 18893
rect 6641 18853 6653 18887
rect 6687 18884 6699 18887
rect 9398 18884 9404 18896
rect 6687 18856 9404 18884
rect 6687 18853 6699 18856
rect 6641 18847 6699 18853
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18785 5687 18819
rect 5629 18779 5687 18785
rect 5644 18680 5672 18779
rect 5718 18776 5724 18828
rect 5776 18816 5782 18828
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5776 18788 5825 18816
rect 5776 18776 5782 18788
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18748 5963 18751
rect 6656 18748 6684 18847
rect 9398 18844 9404 18856
rect 9456 18844 9462 18896
rect 17773 18887 17831 18893
rect 17773 18853 17785 18887
rect 17819 18884 17831 18887
rect 18874 18884 18880 18896
rect 17819 18856 18880 18884
rect 17819 18853 17831 18856
rect 17773 18847 17831 18853
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 7466 18816 7472 18828
rect 7427 18788 7472 18816
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18785 7711 18819
rect 18690 18816 18696 18828
rect 7653 18779 7711 18785
rect 11624 18788 12434 18816
rect 5951 18720 6684 18748
rect 7668 18748 7696 18779
rect 11624 18748 11652 18788
rect 7668 18720 11652 18748
rect 11701 18751 11759 18757
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 11701 18717 11713 18751
rect 11747 18748 11759 18751
rect 12406 18748 12434 18788
rect 17144 18788 18696 18816
rect 13814 18748 13820 18760
rect 11747 18720 11928 18748
rect 12406 18720 13820 18748
rect 11747 18717 11759 18720
rect 11701 18711 11759 18717
rect 10962 18680 10968 18692
rect 5644 18652 10968 18680
rect 7377 18615 7435 18621
rect 7377 18581 7389 18615
rect 7423 18612 7435 18615
rect 7834 18612 7840 18624
rect 7423 18584 7840 18612
rect 7423 18581 7435 18584
rect 7377 18575 7435 18581
rect 7834 18572 7840 18584
rect 7892 18612 7898 18624
rect 8021 18615 8079 18621
rect 8021 18612 8033 18615
rect 7892 18584 8033 18612
rect 7892 18572 7898 18584
rect 8021 18581 8033 18584
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 10336 18621 10364 18652
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 11238 18640 11244 18692
rect 11296 18680 11302 18692
rect 11434 18683 11492 18689
rect 11434 18680 11446 18683
rect 11296 18652 11446 18680
rect 11296 18640 11302 18652
rect 11434 18649 11446 18652
rect 11480 18649 11492 18683
rect 11434 18643 11492 18649
rect 11900 18624 11928 18720
rect 13814 18708 13820 18720
rect 13872 18708 13878 18760
rect 17144 18757 17172 18788
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 19794 18816 19800 18828
rect 19755 18788 19800 18816
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17460 18720 17601 18748
rect 17460 18708 17466 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 17589 18711 17647 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18748 19579 18751
rect 19567 18720 20300 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 18616 18680 18644 18711
rect 20272 18692 20300 18720
rect 20042 18683 20100 18689
rect 20042 18680 20054 18683
rect 17328 18652 18644 18680
rect 18708 18652 20054 18680
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9456 18584 9689 18612
rect 9456 18572 9462 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9677 18575 9735 18581
rect 10321 18615 10379 18621
rect 10321 18581 10333 18615
rect 10367 18581 10379 18615
rect 10321 18575 10379 18581
rect 11882 18572 11888 18624
rect 11940 18612 11946 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11940 18584 11989 18612
rect 11940 18572 11946 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 13170 18612 13176 18624
rect 12124 18584 13176 18612
rect 12124 18572 12130 18584
rect 13170 18572 13176 18584
rect 13228 18612 13234 18624
rect 13538 18612 13544 18624
rect 13228 18584 13544 18612
rect 13228 18572 13234 18584
rect 13538 18572 13544 18584
rect 13596 18612 13602 18624
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 13596 18584 13645 18612
rect 13596 18572 13602 18584
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 16485 18615 16543 18621
rect 16485 18581 16497 18615
rect 16531 18612 16543 18615
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16531 18584 16865 18612
rect 16531 18581 16543 18584
rect 16485 18575 16543 18581
rect 16853 18581 16865 18584
rect 16899 18612 16911 18615
rect 16942 18612 16948 18624
rect 16899 18584 16948 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17328 18621 17356 18652
rect 17313 18615 17371 18621
rect 17313 18581 17325 18615
rect 17359 18581 17371 18615
rect 17313 18575 17371 18581
rect 17862 18572 17868 18624
rect 17920 18612 17926 18624
rect 18708 18612 18736 18652
rect 20042 18649 20054 18652
rect 20088 18649 20100 18683
rect 20042 18643 20100 18649
rect 20254 18640 20260 18692
rect 20312 18640 20318 18692
rect 21542 18680 21548 18692
rect 20364 18652 21548 18680
rect 17920 18584 18736 18612
rect 18785 18615 18843 18621
rect 17920 18572 17926 18584
rect 18785 18581 18797 18615
rect 18831 18612 18843 18615
rect 20364 18612 20392 18652
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 18831 18584 20392 18612
rect 18831 18581 18843 18584
rect 18785 18575 18843 18581
rect 21082 18572 21088 18624
rect 21140 18612 21146 18624
rect 21177 18615 21235 18621
rect 21177 18612 21189 18615
rect 21140 18584 21189 18612
rect 21140 18572 21146 18584
rect 21177 18581 21189 18584
rect 21223 18612 21235 18615
rect 21358 18612 21364 18624
rect 21223 18584 21364 18612
rect 21223 18581 21235 18584
rect 21177 18575 21235 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 7469 18411 7527 18417
rect 7469 18377 7481 18411
rect 7515 18408 7527 18411
rect 7558 18408 7564 18420
rect 7515 18380 7564 18408
rect 7515 18377 7527 18380
rect 7469 18371 7527 18377
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 8481 18411 8539 18417
rect 8481 18377 8493 18411
rect 8527 18408 8539 18411
rect 10502 18408 10508 18420
rect 8527 18380 10508 18408
rect 8527 18377 8539 18380
rect 8481 18371 8539 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 19613 18411 19671 18417
rect 19613 18408 19625 18411
rect 19024 18380 19625 18408
rect 19024 18368 19030 18380
rect 19613 18377 19625 18380
rect 19659 18377 19671 18411
rect 19613 18371 19671 18377
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 6733 18343 6791 18349
rect 6733 18340 6745 18343
rect 6696 18312 6745 18340
rect 6696 18300 6702 18312
rect 6733 18309 6745 18312
rect 6779 18309 6791 18343
rect 10904 18343 10962 18349
rect 10904 18340 10916 18343
rect 6733 18303 6791 18309
rect 8680 18312 10916 18340
rect 8202 18272 8208 18284
rect 6472 18244 8208 18272
rect 5166 18204 5172 18216
rect 5127 18176 5172 18204
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 6472 18213 6500 18244
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18241 8447 18275
rect 8389 18235 8447 18241
rect 6457 18207 6515 18213
rect 6457 18173 6469 18207
rect 6503 18173 6515 18207
rect 6457 18167 6515 18173
rect 6546 18164 6552 18216
rect 6604 18204 6610 18216
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6604 18176 6653 18204
rect 6604 18164 6610 18176
rect 6641 18173 6653 18176
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 8404 18148 8432 18235
rect 8680 18213 8708 18312
rect 10904 18309 10916 18312
rect 10950 18340 10962 18343
rect 11790 18340 11796 18352
rect 10950 18312 11796 18340
rect 10950 18309 10962 18312
rect 10904 18303 10962 18309
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 12710 18300 12716 18352
rect 12768 18340 12774 18352
rect 13050 18343 13108 18349
rect 13050 18340 13062 18343
rect 12768 18312 13062 18340
rect 12768 18300 12774 18312
rect 13050 18309 13062 18312
rect 13096 18309 13108 18343
rect 13050 18303 13108 18309
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 17098 18343 17156 18349
rect 17098 18340 17110 18343
rect 16908 18312 17110 18340
rect 16908 18300 16914 18312
rect 17098 18309 17110 18312
rect 17144 18340 17156 18343
rect 17218 18340 17224 18352
rect 17144 18312 17224 18340
rect 17144 18309 17156 18312
rect 17098 18303 17156 18309
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 9732 18244 11744 18272
rect 9732 18232 9738 18244
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18204 11207 18207
rect 11195 18176 11652 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 5534 18096 5540 18148
rect 5592 18136 5598 18148
rect 8021 18139 8079 18145
rect 8021 18136 8033 18139
rect 5592 18108 8033 18136
rect 5592 18096 5598 18108
rect 8021 18105 8033 18108
rect 8067 18105 8079 18139
rect 8386 18136 8392 18148
rect 8299 18108 8392 18136
rect 8021 18099 8079 18105
rect 8386 18096 8392 18108
rect 8444 18136 8450 18148
rect 9125 18139 9183 18145
rect 9125 18136 9137 18139
rect 8444 18108 9137 18136
rect 8444 18096 8450 18108
rect 9125 18105 9137 18108
rect 9171 18136 9183 18139
rect 9171 18108 9904 18136
rect 9171 18105 9183 18108
rect 9125 18099 9183 18105
rect 7101 18071 7159 18077
rect 7101 18037 7113 18071
rect 7147 18068 7159 18071
rect 8570 18068 8576 18080
rect 7147 18040 8576 18068
rect 7147 18037 7159 18040
rect 7101 18031 7159 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 9766 18068 9772 18080
rect 9727 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 9876 18068 9904 18108
rect 10778 18068 10784 18080
rect 9876 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11624 18077 11652 18176
rect 11716 18136 11744 18244
rect 11882 18232 11888 18284
rect 11940 18272 11946 18284
rect 12805 18275 12863 18281
rect 12805 18272 12817 18275
rect 11940 18244 12817 18272
rect 11940 18232 11946 18244
rect 12805 18241 12817 18244
rect 12851 18241 12863 18275
rect 16942 18272 16948 18284
rect 12805 18235 12863 18241
rect 16868 18244 16948 18272
rect 15930 18204 15936 18216
rect 15891 18176 15936 18204
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 16868 18213 16896 18244
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19024 18244 19165 18272
rect 19024 18232 19030 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19429 18275 19487 18281
rect 19429 18241 19441 18275
rect 19475 18272 19487 18275
rect 19518 18272 19524 18284
rect 19475 18244 19524 18272
rect 19475 18241 19487 18244
rect 19429 18235 19487 18241
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 19760 18244 19993 18272
rect 19760 18232 19766 18244
rect 19981 18241 19993 18244
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 20496 18244 20545 18272
rect 20496 18232 20502 18244
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 21082 18272 21088 18284
rect 21043 18244 21088 18272
rect 20533 18235 20591 18241
rect 21082 18232 21088 18244
rect 21140 18232 21146 18284
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 11716 18108 12434 18136
rect 11609 18071 11667 18077
rect 11609 18037 11621 18071
rect 11655 18068 11667 18071
rect 11882 18068 11888 18080
rect 11655 18040 11888 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 12406 18068 12434 18108
rect 14185 18071 14243 18077
rect 14185 18068 14197 18071
rect 12406 18040 14197 18068
rect 14185 18037 14197 18040
rect 14231 18068 14243 18071
rect 14274 18068 14280 18080
rect 14231 18040 14280 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 14461 18071 14519 18077
rect 14461 18068 14473 18071
rect 14424 18040 14473 18068
rect 14424 18028 14430 18040
rect 14461 18037 14473 18040
rect 14507 18037 14519 18071
rect 16868 18068 16896 18167
rect 18601 18139 18659 18145
rect 18601 18136 18613 18139
rect 17788 18108 18613 18136
rect 17788 18068 17816 18108
rect 18601 18105 18613 18108
rect 18647 18136 18659 18139
rect 19794 18136 19800 18148
rect 18647 18108 19800 18136
rect 18647 18105 18659 18108
rect 18601 18099 18659 18105
rect 19794 18096 19800 18108
rect 19852 18096 19858 18148
rect 20162 18136 20168 18148
rect 20123 18108 20168 18136
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 22462 18136 22468 18148
rect 20548 18108 22468 18136
rect 16868 18040 17816 18068
rect 14461 18031 14519 18037
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18233 18071 18291 18077
rect 18233 18068 18245 18071
rect 17920 18040 18245 18068
rect 17920 18028 17926 18040
rect 18233 18037 18245 18040
rect 18279 18037 18291 18071
rect 18233 18031 18291 18037
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 20548 18068 20576 18108
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 19015 18040 20576 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 20622 18028 20628 18080
rect 20680 18068 20686 18080
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20680 18040 20729 18068
rect 20680 18028 20686 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 21266 18068 21272 18080
rect 21227 18040 21272 18068
rect 20717 18031 20775 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4764 17836 4813 17864
rect 4764 17824 4770 17836
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 9766 17864 9772 17876
rect 4801 17827 4859 17833
rect 5460 17836 9772 17864
rect 5460 17737 5488 17836
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16209 17867 16267 17873
rect 16209 17864 16221 17867
rect 16172 17836 16221 17864
rect 16172 17824 16178 17836
rect 16209 17833 16221 17836
rect 16255 17833 16267 17867
rect 16209 17827 16267 17833
rect 16390 17824 16396 17876
rect 16448 17864 16454 17876
rect 17494 17864 17500 17876
rect 16448 17836 17500 17864
rect 16448 17824 16454 17836
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 18012 17836 19717 17864
rect 18012 17824 18018 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 16850 17796 16856 17808
rect 7392 17768 16856 17796
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 1688 17700 5457 17728
rect 1688 17669 1716 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 6638 17728 6644 17740
rect 6599 17700 6644 17728
rect 5445 17691 5503 17697
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 7392 17737 7420 17768
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 7377 17731 7435 17737
rect 7377 17697 7389 17731
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17728 7527 17731
rect 7742 17728 7748 17740
rect 7515 17700 7748 17728
rect 7515 17697 7527 17700
rect 7469 17691 7527 17697
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 8297 17731 8355 17737
rect 8297 17728 8309 17731
rect 7852 17700 8309 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 1673 17623 1731 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5261 17595 5319 17601
rect 5261 17561 5273 17595
rect 5307 17592 5319 17595
rect 5534 17592 5540 17604
rect 5307 17564 5540 17592
rect 5307 17561 5319 17564
rect 5261 17555 5319 17561
rect 5534 17552 5540 17564
rect 5592 17552 5598 17604
rect 7561 17595 7619 17601
rect 7561 17561 7573 17595
rect 7607 17592 7619 17595
rect 7852 17592 7880 17700
rect 8297 17697 8309 17700
rect 8343 17728 8355 17731
rect 9122 17728 9128 17740
rect 8343 17700 9128 17728
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 17862 17728 17868 17740
rect 15703 17700 17868 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18877 17731 18935 17737
rect 18877 17697 18889 17731
rect 18923 17728 18935 17731
rect 19334 17728 19340 17740
rect 18923 17700 19340 17728
rect 18923 17697 18935 17700
rect 18877 17691 18935 17697
rect 19334 17688 19340 17700
rect 19392 17728 19398 17740
rect 19392 17700 19840 17728
rect 19392 17688 19398 17700
rect 19812 17672 19840 17700
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17660 15899 17663
rect 15930 17660 15936 17672
rect 15887 17632 15936 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 16853 17663 16911 17669
rect 16853 17629 16865 17663
rect 16899 17629 16911 17663
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 16853 17623 16911 17629
rect 17052 17632 19257 17660
rect 15749 17595 15807 17601
rect 15749 17592 15761 17595
rect 7607 17564 7880 17592
rect 7944 17564 15761 17592
rect 7607 17561 7619 17564
rect 7561 17555 7619 17561
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 7944 17533 7972 17564
rect 15749 17561 15761 17564
rect 15795 17561 15807 17595
rect 15749 17555 15807 17561
rect 7929 17527 7987 17533
rect 7929 17493 7941 17527
rect 7975 17493 7987 17527
rect 7929 17487 7987 17493
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 16868 17524 16896 17623
rect 17052 17533 17080 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19794 17620 19800 17672
rect 19852 17660 19858 17672
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 19852 17632 21097 17660
rect 19852 17620 19858 17632
rect 20640 17604 20668 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 18598 17552 18604 17604
rect 18656 17601 18662 17604
rect 18656 17592 18668 17601
rect 18656 17564 18701 17592
rect 18800 17564 20576 17592
rect 18656 17555 18668 17564
rect 18656 17552 18662 17555
rect 8628 17496 16896 17524
rect 17037 17527 17095 17533
rect 8628 17484 8634 17496
rect 17037 17493 17049 17527
rect 17083 17493 17095 17527
rect 17037 17487 17095 17493
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 18800 17524 18828 17564
rect 17552 17496 18828 17524
rect 19429 17527 19487 17533
rect 17552 17484 17558 17496
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19610 17524 19616 17536
rect 19475 17496 19616 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 20548 17524 20576 17564
rect 20622 17552 20628 17604
rect 20680 17552 20686 17604
rect 20818 17595 20876 17601
rect 20818 17592 20830 17595
rect 20732 17564 20830 17592
rect 20732 17524 20760 17564
rect 20818 17561 20830 17564
rect 20864 17561 20876 17595
rect 20818 17555 20876 17561
rect 20548 17496 20760 17524
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 5534 17320 5540 17332
rect 5447 17292 5540 17320
rect 5534 17280 5540 17292
rect 5592 17320 5598 17332
rect 8386 17320 8392 17332
rect 5592 17292 8392 17320
rect 5592 17280 5598 17292
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 16022 17320 16028 17332
rect 15983 17292 16028 17320
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 16761 17323 16819 17329
rect 16761 17289 16773 17323
rect 16807 17320 16819 17323
rect 16942 17320 16948 17332
rect 16807 17292 16948 17320
rect 16807 17289 16819 17292
rect 16761 17283 16819 17289
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 18785 17323 18843 17329
rect 18785 17289 18797 17323
rect 18831 17320 18843 17323
rect 19334 17320 19340 17332
rect 18831 17292 19340 17320
rect 18831 17289 18843 17292
rect 18785 17283 18843 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 19705 17323 19763 17329
rect 19705 17289 19717 17323
rect 19751 17320 19763 17323
rect 21082 17320 21088 17332
rect 19751 17292 21088 17320
rect 19751 17289 19763 17292
rect 19705 17283 19763 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 4798 17212 4804 17264
rect 4856 17252 4862 17264
rect 14124 17255 14182 17261
rect 4856 17224 12434 17252
rect 4856 17212 4862 17224
rect 10870 17144 10876 17196
rect 10928 17193 10934 17196
rect 10928 17184 10940 17193
rect 10928 17156 10973 17184
rect 10928 17147 10940 17156
rect 10928 17144 10934 17147
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11195 17088 11652 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 4154 17008 4160 17060
rect 4212 17048 4218 17060
rect 8018 17048 8024 17060
rect 4212 17020 8024 17048
rect 4212 17008 4218 17020
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 11624 16989 11652 17088
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11882 16980 11888 16992
rect 11655 16952 11888 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12406 16980 12434 17224
rect 14124 17221 14136 17255
rect 14170 17252 14182 17255
rect 14274 17252 14280 17264
rect 14170 17224 14280 17252
rect 14170 17221 14182 17224
rect 14124 17215 14182 17221
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14901 17187 14959 17193
rect 14901 17184 14913 17187
rect 13872 17156 14913 17184
rect 13872 17144 13878 17156
rect 14901 17153 14913 17156
rect 14947 17153 14959 17187
rect 14901 17147 14959 17153
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 15896 17156 19257 17184
rect 15896 17144 15902 17156
rect 19245 17153 19257 17156
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 14366 17116 14372 17128
rect 14327 17088 14372 17116
rect 14366 17076 14372 17088
rect 14424 17116 14430 17128
rect 14645 17119 14703 17125
rect 14645 17116 14657 17119
rect 14424 17088 14657 17116
rect 14424 17076 14430 17088
rect 14645 17085 14657 17088
rect 14691 17085 14703 17119
rect 14645 17079 14703 17085
rect 17678 17008 17684 17060
rect 17736 17048 17742 17060
rect 19061 17051 19119 17057
rect 19061 17048 19073 17051
rect 17736 17020 19073 17048
rect 17736 17008 17742 17020
rect 19061 17017 19073 17020
rect 19107 17017 19119 17051
rect 19061 17011 19119 17017
rect 19536 16992 19564 17147
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19668 17156 19993 17184
rect 19668 17144 19674 17156
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20533 17187 20591 17193
rect 20533 17184 20545 17187
rect 20128 17156 20545 17184
rect 20128 17144 20134 17156
rect 20533 17153 20545 17156
rect 20579 17153 20591 17187
rect 20533 17147 20591 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 20772 17156 21097 17184
rect 20772 17144 20778 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 12986 16980 12992 16992
rect 12406 16952 12992 16980
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 19518 16940 19524 16992
rect 19576 16940 19582 16992
rect 20162 16980 20168 16992
rect 20123 16952 20168 16980
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 20530 16940 20536 16992
rect 20588 16980 20594 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20588 16952 20729 16980
rect 20588 16940 20594 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 20717 16943 20775 16949
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 4614 16736 4620 16788
rect 4672 16776 4678 16788
rect 4672 16748 6132 16776
rect 4672 16736 4678 16748
rect 5810 16708 5816 16720
rect 4908 16680 5816 16708
rect 4798 16640 4804 16652
rect 4759 16612 4804 16640
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 4908 16581 4936 16680
rect 5810 16668 5816 16680
rect 5868 16668 5874 16720
rect 4893 16575 4951 16581
rect 4893 16541 4905 16575
rect 4939 16541 4951 16575
rect 4893 16535 4951 16541
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16572 5043 16575
rect 5534 16572 5540 16584
rect 5031 16544 5540 16572
rect 5031 16541 5043 16544
rect 4985 16535 5043 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 6104 16581 6132 16748
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 18656 16748 19625 16776
rect 18656 16736 18662 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 20680 16748 21036 16776
rect 20680 16736 20686 16748
rect 9766 16708 9772 16720
rect 6288 16680 9772 16708
rect 6288 16649 6316 16680
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 18782 16708 18788 16720
rect 18743 16680 18788 16708
rect 18782 16668 18788 16680
rect 18840 16668 18846 16720
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 7926 16640 7932 16652
rect 6963 16612 7788 16640
rect 7887 16612 7932 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 6089 16575 6147 16581
rect 6089 16541 6101 16575
rect 6135 16541 6147 16575
rect 7760 16572 7788 16612
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 9784 16640 9812 16668
rect 8036 16612 9720 16640
rect 9784 16612 10180 16640
rect 8036 16572 8064 16612
rect 7760 16544 8064 16572
rect 6089 16535 6147 16541
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 8113 16507 8171 16513
rect 8113 16504 8125 16507
rect 7892 16476 8125 16504
rect 7892 16464 7898 16476
rect 8113 16473 8125 16476
rect 8159 16504 8171 16507
rect 8941 16507 8999 16513
rect 8941 16504 8953 16507
rect 8159 16476 8953 16504
rect 8159 16473 8171 16476
rect 8113 16467 8171 16473
rect 8941 16473 8953 16476
rect 8987 16473 8999 16507
rect 9692 16504 9720 16612
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 9824 16544 10057 16572
rect 9824 16532 9830 16544
rect 10045 16541 10057 16544
rect 10091 16541 10103 16575
rect 10152 16572 10180 16612
rect 14366 16600 14372 16652
rect 14424 16600 14430 16652
rect 21008 16649 21036 16748
rect 20993 16643 21051 16649
rect 20993 16609 21005 16643
rect 21039 16640 21051 16643
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 21039 16612 21281 16640
rect 21039 16609 21051 16612
rect 20993 16603 21051 16609
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 10301 16575 10359 16581
rect 10301 16572 10313 16575
rect 10152 16544 10313 16572
rect 10045 16535 10103 16541
rect 10301 16541 10313 16544
rect 10347 16541 10359 16575
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 10301 16535 10359 16541
rect 11882 16532 11888 16544
rect 11940 16572 11946 16584
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 11940 16544 13553 16572
rect 11940 16532 11946 16544
rect 13541 16541 13553 16544
rect 13587 16572 13599 16575
rect 14384 16572 14412 16600
rect 14461 16575 14519 16581
rect 14461 16572 14473 16575
rect 13587 16544 14473 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 14461 16541 14473 16544
rect 14507 16541 14519 16575
rect 18138 16572 18144 16584
rect 18099 16544 18144 16572
rect 14461 16535 14519 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 20737 16575 20795 16581
rect 20737 16541 20749 16575
rect 20783 16572 20795 16575
rect 21358 16572 21364 16584
rect 20783 16544 21364 16572
rect 20783 16541 20795 16544
rect 20737 16535 20795 16541
rect 11698 16504 11704 16516
rect 9692 16476 11704 16504
rect 8941 16467 8999 16473
rect 11698 16464 11704 16476
rect 11756 16504 11762 16516
rect 12130 16507 12188 16513
rect 12130 16504 12142 16507
rect 11756 16476 12142 16504
rect 11756 16464 11762 16476
rect 12130 16473 12142 16476
rect 12176 16473 12188 16507
rect 12130 16467 12188 16473
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 18616 16504 18644 16535
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 12308 16476 18644 16504
rect 12308 16464 12314 16476
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 5353 16439 5411 16445
rect 5353 16436 5365 16439
rect 5316 16408 5365 16436
rect 5316 16396 5322 16408
rect 5353 16405 5365 16408
rect 5399 16405 5411 16439
rect 5626 16436 5632 16448
rect 5587 16408 5632 16436
rect 5353 16399 5411 16405
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 5994 16436 6000 16448
rect 5955 16408 6000 16436
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 7006 16436 7012 16448
rect 6967 16408 7012 16436
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7101 16439 7159 16445
rect 7101 16405 7113 16439
rect 7147 16436 7159 16439
rect 7282 16436 7288 16448
rect 7147 16408 7288 16436
rect 7147 16405 7159 16408
rect 7101 16399 7159 16405
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 7466 16436 7472 16448
rect 7427 16408 7472 16436
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 8481 16439 8539 16445
rect 8481 16436 8493 16439
rect 8444 16408 8493 16436
rect 8444 16396 8450 16408
rect 8481 16405 8493 16408
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 11296 16408 11437 16436
rect 11296 16396 11302 16408
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 11425 16399 11483 16405
rect 13265 16439 13323 16445
rect 13265 16405 13277 16439
rect 13311 16436 13323 16439
rect 13814 16436 13820 16448
rect 13311 16408 13820 16436
rect 13311 16405 13323 16408
rect 13265 16399 13323 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 18325 16439 18383 16445
rect 18325 16405 18337 16439
rect 18371 16436 18383 16439
rect 19518 16436 19524 16448
rect 18371 16408 19524 16436
rect 18371 16405 18383 16408
rect 18325 16399 18383 16405
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 5258 16232 5264 16244
rect 5219 16204 5264 16232
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 7282 16232 7288 16244
rect 7243 16204 7288 16232
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 8386 16232 8392 16244
rect 8347 16204 8392 16232
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 12250 16232 12256 16244
rect 8895 16204 12256 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 12406 16204 14136 16232
rect 12406 16164 12434 16204
rect 5184 16136 12434 16164
rect 5184 16037 5212 16136
rect 12986 16124 12992 16176
rect 13044 16164 13050 16176
rect 13602 16167 13660 16173
rect 13602 16164 13614 16167
rect 13044 16136 13614 16164
rect 13044 16124 13050 16136
rect 13602 16133 13614 16136
rect 13648 16133 13660 16167
rect 14108 16164 14136 16204
rect 14366 16192 14372 16244
rect 14424 16232 14430 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14424 16204 15025 16232
rect 14424 16192 14430 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 18969 16235 19027 16241
rect 18969 16201 18981 16235
rect 19015 16201 19027 16235
rect 18969 16195 19027 16201
rect 19429 16235 19487 16241
rect 19429 16201 19441 16235
rect 19475 16232 19487 16235
rect 20070 16232 20076 16244
rect 19475 16204 20076 16232
rect 19475 16201 19487 16204
rect 19429 16195 19487 16201
rect 15286 16164 15292 16176
rect 14108 16136 15292 16164
rect 13602 16127 13660 16133
rect 15286 16124 15292 16136
rect 15344 16124 15350 16176
rect 18984 16164 19012 16195
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20257 16235 20315 16241
rect 20257 16201 20269 16235
rect 20303 16232 20315 16235
rect 20622 16232 20628 16244
rect 20303 16204 20628 16232
rect 20303 16201 20315 16204
rect 20257 16195 20315 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20714 16164 20720 16176
rect 18984 16136 20720 16164
rect 20714 16124 20720 16136
rect 20772 16124 20778 16176
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 5442 16096 5448 16108
rect 5399 16068 5448 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 9125 16099 9183 16105
rect 9125 16096 9137 16099
rect 8527 16068 9137 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 9125 16065 9137 16068
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 17497 16099 17555 16105
rect 17497 16065 17509 16099
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 16028 8355 16031
rect 10870 16028 10876 16040
rect 8343 16000 10876 16028
rect 8343 15997 8355 16000
rect 8297 15991 8355 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 13357 16031 13415 16037
rect 13357 16028 13369 16031
rect 11940 16000 13369 16028
rect 11940 15988 11946 16000
rect 13357 15997 13369 16000
rect 13403 15997 13415 16031
rect 13357 15991 13415 15997
rect 5721 15963 5779 15969
rect 5721 15929 5733 15963
rect 5767 15960 5779 15963
rect 17512 15960 17540 16059
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 18012 16068 18153 16096
rect 18012 16056 18018 16068
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18141 16059 18199 16065
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16096 19303 16099
rect 19291 16068 19748 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 19720 15969 19748 16068
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19852 16068 19901 16096
rect 19852 16056 19858 16068
rect 19889 16065 19901 16068
rect 19935 16065 19947 16099
rect 20530 16096 20536 16108
rect 20491 16068 20536 16096
rect 19889 16059 19947 16065
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 20346 15988 20352 16040
rect 20404 16028 20410 16040
rect 21100 16028 21128 16059
rect 20404 16000 21128 16028
rect 20404 15988 20410 16000
rect 5767 15932 12434 15960
rect 5767 15929 5779 15932
rect 5721 15923 5779 15929
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6052 15864 6561 15892
rect 6052 15852 6058 15864
rect 6549 15861 6561 15864
rect 6595 15892 6607 15895
rect 9122 15892 9128 15904
rect 6595 15864 9128 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 11514 15892 11520 15904
rect 11475 15864 11520 15892
rect 11514 15852 11520 15864
rect 11572 15892 11578 15904
rect 11882 15892 11888 15904
rect 11572 15864 11888 15892
rect 11572 15852 11578 15864
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12406 15892 12434 15932
rect 14660 15932 17540 15960
rect 19705 15963 19763 15969
rect 14660 15892 14688 15932
rect 19705 15929 19717 15963
rect 19751 15929 19763 15963
rect 19705 15923 19763 15929
rect 12406 15864 14688 15892
rect 14737 15895 14795 15901
rect 14737 15861 14749 15895
rect 14783 15892 14795 15895
rect 15286 15892 15292 15904
rect 14783 15864 15292 15892
rect 14783 15861 14795 15864
rect 14737 15855 14795 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 17678 15892 17684 15904
rect 17639 15864 17684 15892
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 18230 15852 18236 15904
rect 18288 15892 18294 15904
rect 18325 15895 18383 15901
rect 18325 15892 18337 15895
rect 18288 15864 18337 15892
rect 18288 15852 18294 15864
rect 18325 15861 18337 15864
rect 18371 15861 18383 15895
rect 20714 15892 20720 15904
rect 20675 15864 20720 15892
rect 18325 15855 18383 15861
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7653 15691 7711 15697
rect 7653 15688 7665 15691
rect 7064 15660 7665 15688
rect 7064 15648 7070 15660
rect 7653 15657 7665 15660
rect 7699 15657 7711 15691
rect 12250 15688 12256 15700
rect 7653 15651 7711 15657
rect 8312 15660 12256 15688
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 8312 15561 8340 15660
rect 12250 15648 12256 15660
rect 12308 15688 12314 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 12308 15660 12357 15688
rect 12308 15648 12314 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 18417 15691 18475 15697
rect 18417 15657 18429 15691
rect 18463 15688 18475 15691
rect 19058 15688 19064 15700
rect 18463 15660 19064 15688
rect 18463 15657 18475 15660
rect 18417 15651 18475 15657
rect 19058 15648 19064 15660
rect 19116 15648 19122 15700
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 20533 15691 20591 15697
rect 20533 15688 20545 15691
rect 20496 15660 20545 15688
rect 20496 15648 20502 15660
rect 20533 15657 20545 15660
rect 20579 15657 20591 15691
rect 20533 15651 20591 15657
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 7708 15524 8125 15552
rect 7708 15512 7714 15524
rect 8113 15521 8125 15524
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 17736 15524 20392 15552
rect 17736 15512 17742 15524
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15484 9830 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 9824 15456 11437 15484
rect 9824 15444 9830 15456
rect 11425 15453 11437 15456
rect 11471 15484 11483 15487
rect 11514 15484 11520 15496
rect 11471 15456 11520 15484
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 11514 15444 11520 15456
rect 11572 15484 11578 15496
rect 12342 15484 12348 15496
rect 11572 15456 12348 15484
rect 11572 15444 11578 15456
rect 12342 15444 12348 15456
rect 12400 15484 12406 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 12400 15456 13737 15484
rect 12400 15444 12406 15456
rect 13725 15453 13737 15456
rect 13771 15484 13783 15487
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13771 15456 14105 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 17037 15487 17095 15493
rect 17037 15453 17049 15487
rect 17083 15484 17095 15487
rect 18230 15484 18236 15496
rect 17083 15456 17448 15484
rect 18191 15456 18236 15484
rect 17083 15453 17095 15456
rect 17037 15447 17095 15453
rect 10042 15425 10048 15428
rect 10036 15379 10048 15425
rect 10100 15416 10106 15428
rect 10100 15388 10136 15416
rect 10042 15376 10048 15379
rect 10100 15376 10106 15388
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 13458 15419 13516 15425
rect 13458 15416 13470 15419
rect 12860 15388 13470 15416
rect 12860 15376 12866 15388
rect 13458 15385 13470 15388
rect 13504 15385 13516 15419
rect 13458 15379 13516 15385
rect 16390 15376 16396 15428
rect 16448 15416 16454 15428
rect 16770 15419 16828 15425
rect 16770 15416 16782 15419
rect 16448 15388 16782 15416
rect 16448 15376 16454 15388
rect 16770 15385 16782 15388
rect 16816 15385 16828 15419
rect 16770 15379 16828 15385
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15348 8079 15351
rect 8386 15348 8392 15360
rect 8067 15320 8392 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 8386 15308 8392 15320
rect 8444 15348 8450 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8444 15320 8953 15348
rect 8444 15308 8450 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11149 15351 11207 15357
rect 11149 15348 11161 15351
rect 11112 15320 11161 15348
rect 11112 15308 11118 15320
rect 11149 15317 11161 15320
rect 11195 15317 11207 15351
rect 11149 15311 11207 15317
rect 15657 15351 15715 15357
rect 15657 15317 15669 15351
rect 15703 15348 15715 15351
rect 15838 15348 15844 15360
rect 15703 15320 15844 15348
rect 15703 15317 15715 15320
rect 15657 15311 15715 15317
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 17420 15357 17448 15456
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 20364 15493 20392 15524
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 22186 15484 22192 15496
rect 21131 15456 22192 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 20088 15416 20116 15447
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 20714 15416 20720 15428
rect 20088 15388 20720 15416
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 17405 15351 17463 15357
rect 17405 15317 17417 15351
rect 17451 15348 17463 15351
rect 17862 15348 17868 15360
rect 17451 15320 17868 15348
rect 17451 15317 17463 15320
rect 17405 15311 17463 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 5537 15147 5595 15153
rect 5537 15113 5549 15147
rect 5583 15144 5595 15147
rect 5626 15144 5632 15156
rect 5583 15116 5632 15144
rect 5583 15113 5595 15116
rect 5537 15107 5595 15113
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 17126 15144 17132 15156
rect 6043 15116 16160 15144
rect 17087 15116 17132 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 7926 15036 7932 15088
rect 7984 15076 7990 15088
rect 9582 15076 9588 15088
rect 7984 15048 9588 15076
rect 7984 15036 7990 15048
rect 9582 15036 9588 15048
rect 9640 15076 9646 15088
rect 9922 15079 9980 15085
rect 9922 15076 9934 15079
rect 9640 15048 9934 15076
rect 9640 15036 9646 15048
rect 9922 15045 9934 15048
rect 9968 15045 9980 15079
rect 9922 15039 9980 15045
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 12400 15048 12940 15076
rect 12400 15036 12406 15048
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5675 14980 6377 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 9766 15008 9772 15020
rect 9723 14980 9772 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12630 15011 12688 15017
rect 12630 15008 12642 15011
rect 12308 14980 12642 15008
rect 12308 14968 12314 14980
rect 12630 14977 12642 14980
rect 12676 14977 12688 15011
rect 12630 14971 12688 14977
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5491 14912 7052 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 7024 14804 7052 14912
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 12912 14949 12940 15048
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 7156 14912 7205 14940
rect 7156 14900 7162 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14940 12955 14943
rect 12943 14912 13308 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 11057 14875 11115 14881
rect 11057 14872 11069 14875
rect 10928 14844 11069 14872
rect 10928 14832 10934 14844
rect 11057 14841 11069 14844
rect 11103 14841 11115 14875
rect 11057 14835 11115 14841
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14872 11575 14875
rect 11698 14872 11704 14884
rect 11563 14844 11704 14872
rect 11563 14841 11575 14844
rect 11517 14835 11575 14841
rect 11698 14832 11704 14844
rect 11756 14832 11762 14884
rect 11238 14804 11244 14816
rect 7024 14776 11244 14804
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 13280 14813 13308 14912
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 14274 14804 14280 14816
rect 13311 14776 14280 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 16132 14804 16160 15116
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 20162 15144 20168 15156
rect 17236 15116 20168 15144
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 17236 15008 17264 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20530 15144 20536 15156
rect 20491 15116 20536 15144
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 17236 14980 17325 15008
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 17552 14980 20085 15008
rect 17552 14968 17558 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 22094 15008 22100 15020
rect 21131 14980 22100 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 20732 14940 20760 14971
rect 22094 14968 22100 14980
rect 22152 14968 22158 15020
rect 16868 14912 20760 14940
rect 16868 14881 16896 14912
rect 16853 14875 16911 14881
rect 16853 14841 16865 14875
rect 16899 14841 16911 14875
rect 16853 14835 16911 14841
rect 20257 14875 20315 14881
rect 20257 14841 20269 14875
rect 20303 14872 20315 14875
rect 20806 14872 20812 14884
rect 20303 14844 20812 14872
rect 20303 14841 20315 14844
rect 20257 14835 20315 14841
rect 20806 14832 20812 14844
rect 20864 14832 20870 14884
rect 19794 14804 19800 14816
rect 16132 14776 19800 14804
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 7837 14603 7895 14609
rect 7837 14569 7849 14603
rect 7883 14600 7895 14603
rect 16666 14600 16672 14612
rect 7883 14572 16672 14600
rect 7883 14569 7895 14572
rect 7837 14563 7895 14569
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 17494 14600 17500 14612
rect 16899 14572 17500 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19518 14600 19524 14612
rect 19383 14572 19524 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19518 14560 19524 14572
rect 19576 14600 19582 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 19576 14572 20269 14600
rect 19576 14560 19582 14572
rect 20257 14569 20269 14572
rect 20303 14600 20315 14603
rect 20622 14600 20628 14612
rect 20303 14572 20628 14600
rect 20303 14569 20315 14572
rect 20257 14563 20315 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 11054 14464 11060 14476
rect 7331 14436 11060 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16393 14467 16451 14473
rect 16393 14464 16405 14467
rect 16071 14436 16405 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16393 14433 16405 14436
rect 16439 14464 16451 14467
rect 16439 14436 17356 14464
rect 16439 14433 16451 14436
rect 16393 14427 16451 14433
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 17328 14405 17356 14436
rect 15758 14399 15816 14405
rect 7616 14368 14780 14396
rect 7616 14356 7622 14368
rect 7469 14331 7527 14337
rect 7469 14297 7481 14331
rect 7515 14328 7527 14331
rect 8113 14331 8171 14337
rect 8113 14328 8125 14331
rect 7515 14300 8125 14328
rect 7515 14297 7527 14300
rect 7469 14291 7527 14297
rect 8113 14297 8125 14300
rect 8159 14297 8171 14331
rect 8113 14291 8171 14297
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 11238 14260 11244 14272
rect 11199 14232 11244 14260
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 14642 14260 14648 14272
rect 14603 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 14752 14260 14780 14368
rect 15758 14365 15770 14399
rect 15804 14365 15816 14399
rect 15758 14359 15816 14365
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 17313 14399 17371 14405
rect 17313 14365 17325 14399
rect 17359 14396 17371 14399
rect 17862 14396 17868 14408
rect 17359 14368 17868 14396
rect 17359 14365 17371 14368
rect 17313 14359 17371 14365
rect 15764 14328 15792 14359
rect 15838 14328 15844 14340
rect 15764 14300 15844 14328
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 16684 14260 16712 14359
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20128 14368 20821 14396
rect 20128 14356 20134 14368
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14396 21143 14399
rect 21634 14396 21640 14408
rect 21131 14368 21640 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 17034 14288 17040 14340
rect 17092 14328 17098 14340
rect 17558 14331 17616 14337
rect 17558 14328 17570 14331
rect 17092 14300 17570 14328
rect 17092 14288 17098 14300
rect 17558 14297 17570 14300
rect 17604 14297 17616 14331
rect 17558 14291 17616 14297
rect 14752 14232 16712 14260
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 18782 14260 18788 14272
rect 18739 14232 18788 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19610 14220 19616 14272
rect 19668 14260 19674 14272
rect 20625 14263 20683 14269
rect 20625 14260 20637 14263
rect 19668 14232 20637 14260
rect 19668 14220 19674 14232
rect 20625 14229 20637 14232
rect 20671 14229 20683 14263
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 20625 14223 20683 14229
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 7098 14056 7104 14068
rect 7059 14028 7104 14056
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7558 14056 7564 14068
rect 7515 14028 7564 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 8294 14056 8300 14068
rect 8255 14028 8300 14056
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 9582 14056 9588 14068
rect 9543 14028 9588 14056
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11296 14028 11529 14056
rect 11296 14016 11302 14028
rect 11517 14025 11529 14028
rect 11563 14056 11575 14059
rect 11606 14056 11612 14068
rect 11563 14028 11612 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12802 14056 12808 14068
rect 12763 14028 12808 14056
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 19245 14059 19303 14065
rect 19245 14025 19257 14059
rect 19291 14056 19303 14059
rect 19291 14028 20024 14056
rect 19291 14025 19303 14028
rect 19245 14019 19303 14025
rect 10720 13991 10778 13997
rect 10720 13957 10732 13991
rect 10766 13988 10778 13991
rect 11054 13988 11060 14000
rect 10766 13960 11060 13988
rect 10766 13957 10778 13960
rect 10720 13951 10778 13957
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 8110 13920 8116 13932
rect 8071 13892 8116 13920
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11256 13920 11284 14016
rect 11790 13948 11796 14000
rect 11848 13988 11854 14000
rect 13940 13991 13998 13997
rect 13940 13988 13952 13991
rect 11848 13960 13952 13988
rect 11848 13948 11854 13960
rect 13940 13957 13952 13960
rect 13986 13988 13998 13991
rect 14642 13988 14648 14000
rect 13986 13960 14648 13988
rect 13986 13957 13998 13960
rect 13940 13951 13998 13957
rect 14642 13948 14648 13960
rect 14700 13948 14706 14000
rect 18132 13991 18190 13997
rect 18132 13957 18144 13991
rect 18178 13988 18190 13991
rect 19886 13988 19892 14000
rect 18178 13960 19892 13988
rect 18178 13957 18190 13960
rect 18132 13951 18190 13957
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 19518 13920 19524 13932
rect 11011 13892 11284 13920
rect 19479 13892 19524 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 19788 13923 19846 13929
rect 19788 13889 19800 13923
rect 19834 13920 19846 13923
rect 19996 13920 20024 14028
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20864 14028 20913 14056
rect 20864 14016 20870 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 21174 14056 21180 14068
rect 21135 14028 21180 14056
rect 20901 14019 20959 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 20622 13920 20628 13932
rect 19834 13892 20628 13920
rect 19834 13889 19846 13892
rect 19788 13883 19846 13889
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 21450 13920 21456 13932
rect 21407 13892 21456 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 6825 13815 6883 13821
rect 6840 13784 6868 13815
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13852 14243 13855
rect 14274 13852 14280 13864
rect 14231 13824 14280 13852
rect 14231 13821 14243 13824
rect 14185 13815 14243 13821
rect 14274 13812 14280 13824
rect 14332 13852 14338 13864
rect 16761 13855 16819 13861
rect 14332 13824 14596 13852
rect 14332 13812 14338 13824
rect 12802 13784 12808 13796
rect 6840 13756 9720 13784
rect 9692 13716 9720 13756
rect 12406 13756 12808 13784
rect 12406 13716 12434 13756
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 14568 13725 14596 13824
rect 16761 13821 16773 13855
rect 16807 13852 16819 13855
rect 17862 13852 17868 13864
rect 16807 13824 17868 13852
rect 16807 13821 16819 13824
rect 16761 13815 16819 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 9692 13688 12434 13716
rect 14553 13719 14611 13725
rect 14553 13685 14565 13719
rect 14599 13716 14611 13719
rect 15010 13716 15016 13728
rect 14599 13688 15016 13716
rect 14599 13685 14611 13688
rect 14553 13679 14611 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7432 13484 7665 13512
rect 7432 13472 7438 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 7653 13475 7711 13481
rect 8220 13484 9965 13512
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 8220 13385 8248 13484
rect 9953 13481 9965 13484
rect 9999 13512 10011 13515
rect 10042 13512 10048 13524
rect 9999 13484 10048 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 11606 13512 11612 13524
rect 11567 13484 11612 13512
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13512 13507 13515
rect 16390 13512 16396 13524
rect 13495 13484 15976 13512
rect 16351 13484 16396 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 4028 13348 8125 13376
rect 4028 13336 4034 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13345 8263 13379
rect 8205 13339 8263 13345
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11624 13376 11652 13472
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11379 13348 12081 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 8021 13243 8079 13249
rect 8021 13209 8033 13243
rect 8067 13240 8079 13243
rect 8386 13240 8392 13252
rect 8067 13212 8392 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 8386 13200 8392 13212
rect 8444 13240 8450 13252
rect 8444 13212 9076 13240
rect 8444 13200 8450 13212
rect 9048 13181 9076 13212
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 11066 13243 11124 13249
rect 11066 13240 11078 13243
rect 9824 13212 11078 13240
rect 9824 13200 9830 13212
rect 11066 13209 11078 13212
rect 11112 13209 11124 13243
rect 11066 13203 11124 13209
rect 11882 13200 11888 13252
rect 11940 13240 11946 13252
rect 12314 13243 12372 13249
rect 12314 13240 12326 13243
rect 11940 13212 12326 13240
rect 11940 13200 11946 13212
rect 12314 13209 12326 13212
rect 12360 13209 12372 13243
rect 12314 13203 12372 13209
rect 9033 13175 9091 13181
rect 9033 13141 9045 13175
rect 9079 13172 9091 13175
rect 11974 13172 11980 13184
rect 9079 13144 11980 13172
rect 9079 13141 9091 13144
rect 9033 13135 9091 13141
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 13464 13172 13492 13475
rect 15948 13444 15976 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 18877 13515 18935 13521
rect 17920 13484 18092 13512
rect 17920 13472 17926 13484
rect 17034 13444 17040 13456
rect 15948 13416 17040 13444
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 18064 13385 18092 13484
rect 18877 13481 18889 13515
rect 18923 13512 18935 13515
rect 19337 13515 19395 13521
rect 19337 13512 19349 13515
rect 18923 13484 19349 13512
rect 18923 13481 18935 13484
rect 18877 13475 18935 13481
rect 19337 13481 19349 13484
rect 19383 13512 19395 13515
rect 19518 13512 19524 13524
rect 19383 13484 19524 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 18892 13376 18920 13475
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 20254 13472 20260 13524
rect 20312 13512 20318 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 20312 13484 20637 13512
rect 20312 13472 20318 13484
rect 20625 13481 20637 13484
rect 20671 13481 20683 13515
rect 21266 13512 21272 13524
rect 21227 13484 21272 13512
rect 20625 13475 20683 13481
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 18095 13348 18920 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 14185 13311 14243 13317
rect 14185 13277 14197 13311
rect 14231 13308 14243 13311
rect 15010 13308 15016 13320
rect 14231 13280 15016 13308
rect 14231 13277 14243 13280
rect 14185 13271 14243 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 15286 13317 15292 13320
rect 15280 13271 15292 13317
rect 15344 13308 15350 13320
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 15344 13280 15380 13308
rect 18064 13280 18521 13308
rect 15286 13268 15292 13271
rect 15344 13268 15350 13280
rect 18064 13252 18092 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 20346 13308 20352 13320
rect 19935 13280 20352 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20346 13268 20352 13280
rect 20404 13268 20410 13320
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 20990 13308 20996 13320
rect 20855 13280 20996 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 21174 13308 21180 13320
rect 21131 13280 21180 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 14826 13200 14832 13252
rect 14884 13240 14890 13252
rect 14884 13212 16804 13240
rect 14884 13200 14890 13212
rect 12124 13144 13492 13172
rect 12124 13132 12130 13144
rect 16482 13132 16488 13184
rect 16540 13172 16546 13184
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 16540 13144 16681 13172
rect 16540 13132 16546 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 16776 13172 16804 13212
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17782 13243 17840 13249
rect 17782 13240 17794 13243
rect 17092 13212 17794 13240
rect 17092 13200 17098 13212
rect 17782 13209 17794 13212
rect 17828 13209 17840 13243
rect 17782 13203 17840 13209
rect 18046 13200 18052 13252
rect 18104 13200 18110 13252
rect 18325 13175 18383 13181
rect 18325 13172 18337 13175
rect 16776 13144 18337 13172
rect 16669 13135 16727 13141
rect 18325 13141 18337 13144
rect 18371 13141 18383 13175
rect 18325 13135 18383 13141
rect 18690 13132 18696 13184
rect 18748 13172 18754 13184
rect 20165 13175 20223 13181
rect 20165 13172 20177 13175
rect 18748 13144 20177 13172
rect 18748 13132 18754 13144
rect 20165 13141 20177 13144
rect 20211 13141 20223 13175
rect 20165 13135 20223 13141
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 7064 12940 7205 12968
rect 7064 12928 7070 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7340 12940 7665 12968
rect 7340 12928 7346 12940
rect 7653 12937 7665 12940
rect 7699 12937 7711 12971
rect 7653 12931 7711 12937
rect 11609 12971 11667 12977
rect 11609 12937 11621 12971
rect 11655 12968 11667 12971
rect 11698 12968 11704 12980
rect 11655 12940 11704 12968
rect 11655 12937 11667 12940
rect 11609 12931 11667 12937
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 8018 12832 8024 12844
rect 7607 12804 8024 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 8018 12792 8024 12804
rect 8076 12832 8082 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8076 12804 8677 12832
rect 8076 12792 8082 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10882 12835 10940 12841
rect 10882 12832 10894 12835
rect 10192 12804 10894 12832
rect 10192 12792 10198 12804
rect 10882 12801 10894 12804
rect 10928 12832 10940 12835
rect 11149 12835 11207 12841
rect 10928 12804 11100 12832
rect 10928 12801 10940 12804
rect 10882 12795 10940 12801
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 8202 12764 8208 12776
rect 8163 12736 8208 12764
rect 7837 12727 7895 12733
rect 7852 12696 7880 12727
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 11072 12764 11100 12804
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11624 12832 11652 12931
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 13814 12968 13820 12980
rect 12032 12940 13820 12968
rect 12032 12928 12038 12940
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 16390 12968 16396 12980
rect 13924 12940 16396 12968
rect 13924 12900 13952 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 18509 12971 18567 12977
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 19518 12968 19524 12980
rect 18555 12940 19524 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 15010 12900 15016 12912
rect 11195 12804 11652 12832
rect 12406 12872 13952 12900
rect 14016 12872 15016 12900
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 12406 12764 12434 12872
rect 14016 12841 14044 12872
rect 15010 12860 15016 12872
rect 15068 12900 15074 12912
rect 15749 12903 15807 12909
rect 15749 12900 15761 12903
rect 15068 12872 15761 12900
rect 15068 12860 15074 12872
rect 15749 12869 15761 12872
rect 15795 12900 15807 12903
rect 18524 12900 18552 12931
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 20036 12940 20085 12968
rect 20036 12928 20042 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 20717 12971 20775 12977
rect 20717 12937 20729 12971
rect 20763 12968 20775 12971
rect 21082 12968 21088 12980
rect 20763 12940 21088 12968
rect 20763 12937 20775 12940
rect 20717 12931 20775 12937
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 15795 12872 18552 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 14274 12841 14280 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14268 12795 14280 12841
rect 14332 12832 14338 12844
rect 16776 12841 16804 12872
rect 16761 12835 16819 12841
rect 14332 12804 14368 12832
rect 14274 12792 14280 12795
rect 14332 12792 14338 12804
rect 16761 12801 16773 12835
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 17028 12835 17086 12841
rect 17028 12801 17040 12835
rect 17074 12832 17086 12835
rect 18782 12832 18788 12844
rect 17074 12804 18788 12832
rect 17074 12801 17086 12804
rect 17028 12795 17086 12801
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 20530 12832 20536 12844
rect 20491 12804 20536 12832
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 21082 12832 21088 12844
rect 21043 12804 21088 12832
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 11072 12736 12434 12764
rect 7852 12668 9904 12696
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 9766 12628 9772 12640
rect 5592 12600 9772 12628
rect 5592 12588 5598 12600
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 9876 12628 9904 12668
rect 11790 12628 11796 12640
rect 9876 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14918 12628 14924 12640
rect 13872 12600 14924 12628
rect 13872 12588 13878 12600
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12628 15439 12631
rect 17034 12628 17040 12640
rect 15427 12600 17040 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 18141 12631 18199 12637
rect 18141 12597 18153 12631
rect 18187 12628 18199 12631
rect 18874 12628 18880 12640
rect 18187 12600 18880 12628
rect 18187 12597 18199 12600
rect 18141 12591 18199 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19797 12631 19855 12637
rect 19797 12597 19809 12631
rect 19843 12628 19855 12631
rect 21358 12628 21364 12640
rect 19843 12600 21364 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 21358 12588 21364 12600
rect 21416 12588 21422 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 12066 12424 12072 12436
rect 7668 12396 12072 12424
rect 6380 12328 6914 12356
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 5534 12288 5540 12300
rect 4939 12260 5540 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 6380 12297 6408 12328
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 5960 12260 6193 12288
rect 5960 12248 5966 12260
rect 6181 12257 6193 12260
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6886 12220 6914 12328
rect 7668 12297 7696 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 20254 12424 20260 12436
rect 20215 12396 20260 12424
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 20898 12424 20904 12436
rect 20859 12396 20904 12424
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 21048 12396 21189 12424
rect 21048 12384 21054 12396
rect 21177 12393 21189 12396
rect 21223 12393 21235 12427
rect 21177 12387 21235 12393
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20530 12356 20536 12368
rect 20027 12328 20536 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12257 7711 12291
rect 10134 12288 10140 12300
rect 7653 12251 7711 12257
rect 7760 12260 10140 12288
rect 7760 12220 7788 12260
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 14550 12288 14556 12300
rect 11072 12260 14556 12288
rect 6886 12192 7788 12220
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8202 12220 8208 12232
rect 7883 12192 8208 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 10893 12223 10951 12229
rect 10893 12220 10905 12223
rect 8352 12192 10905 12220
rect 8352 12180 8358 12192
rect 10893 12189 10905 12192
rect 10939 12220 10951 12223
rect 11072 12220 11100 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 10939 12192 11100 12220
rect 11149 12223 11207 12229
rect 10939 12189 10951 12192
rect 10893 12183 10951 12189
rect 11149 12189 11161 12223
rect 11195 12220 11207 12223
rect 11195 12192 11560 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 4985 12155 5043 12161
rect 4985 12121 4997 12155
rect 5031 12152 5043 12155
rect 6089 12155 6147 12161
rect 5031 12124 5764 12152
rect 5031 12121 5043 12124
rect 4985 12115 5043 12121
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5442 12084 5448 12096
rect 5132 12056 5177 12084
rect 5403 12056 5448 12084
rect 5132 12044 5138 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5736 12093 5764 12124
rect 6089 12121 6101 12155
rect 6135 12152 6147 12155
rect 6733 12155 6791 12161
rect 6733 12152 6745 12155
rect 6135 12124 6745 12152
rect 6135 12121 6147 12124
rect 6089 12115 6147 12121
rect 6733 12121 6745 12124
rect 6779 12121 6791 12155
rect 6733 12115 6791 12121
rect 7745 12155 7803 12161
rect 7745 12121 7757 12155
rect 7791 12152 7803 12155
rect 10502 12152 10508 12164
rect 7791 12124 10508 12152
rect 7791 12121 7803 12124
rect 7745 12115 7803 12121
rect 5721 12087 5779 12093
rect 5721 12053 5733 12087
rect 5767 12053 5779 12087
rect 6748 12084 6776 12115
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 8018 12084 8024 12096
rect 6748 12056 8024 12084
rect 5721 12047 5779 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 9766 12084 9772 12096
rect 9727 12056 9772 12084
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 11532 12093 11560 12192
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 15010 12220 15016 12232
rect 13964 12192 15016 12220
rect 13964 12180 13970 12192
rect 15010 12180 15016 12192
rect 15068 12220 15074 12232
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 15068 12192 15577 12220
rect 15068 12180 15074 12192
rect 15565 12189 15577 12192
rect 15611 12220 15623 12223
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15611 12192 15853 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 15841 12183 15899 12189
rect 19536 12192 19809 12220
rect 15320 12155 15378 12161
rect 15320 12121 15332 12155
rect 15366 12152 15378 12155
rect 16114 12152 16120 12164
rect 15366 12124 16120 12152
rect 15366 12121 15378 12124
rect 15320 12115 15378 12121
rect 16114 12112 16120 12124
rect 16172 12112 16178 12164
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 11698 12084 11704 12096
rect 11563 12056 11704 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 14185 12087 14243 12093
rect 14185 12053 14197 12087
rect 14231 12084 14243 12087
rect 14274 12084 14280 12096
rect 14231 12056 14280 12084
rect 14231 12053 14243 12056
rect 14185 12047 14243 12053
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 19536 12093 19564 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 21174 12220 21180 12232
rect 20763 12192 21180 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 20456 12152 20484 12183
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 21358 12220 21364 12232
rect 21319 12192 21364 12220
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 21542 12152 21548 12164
rect 20456 12124 21548 12152
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 19116 12056 19533 12084
rect 19116 12044 19122 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 21634 12044 21640 12096
rect 21692 12084 21698 12096
rect 22278 12084 22284 12096
rect 21692 12056 22284 12084
rect 21692 12044 21698 12056
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 5132 11852 5549 11880
rect 5132 11840 5138 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 5537 11843 5595 11849
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8662 11880 8668 11892
rect 7975 11852 8668 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 13906 11880 13912 11892
rect 13867 11852 13912 11880
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 18690 11840 18696 11892
rect 18748 11880 18754 11892
rect 18966 11880 18972 11892
rect 18748 11852 18972 11880
rect 18748 11840 18754 11852
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 21361 11883 21419 11889
rect 21361 11849 21373 11883
rect 21407 11880 21419 11883
rect 21542 11880 21548 11892
rect 21407 11852 21548 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 20806 11821 20812 11824
rect 20748 11815 20812 11821
rect 20748 11781 20760 11815
rect 20794 11781 20812 11815
rect 20748 11775 20812 11781
rect 20806 11772 20812 11775
rect 20864 11772 20870 11824
rect 21266 11772 21272 11824
rect 21324 11812 21330 11824
rect 21634 11812 21640 11824
rect 21324 11784 21640 11812
rect 21324 11772 21330 11784
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8202 11744 8208 11756
rect 7791 11716 8208 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11744 18567 11747
rect 21358 11744 21364 11756
rect 18555 11716 21364 11744
rect 18555 11713 18567 11716
rect 18509 11707 18567 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 20993 11679 21051 11685
rect 20993 11645 21005 11679
rect 21039 11676 21051 11679
rect 21266 11676 21272 11688
rect 21039 11648 21272 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 18782 11540 18788 11552
rect 18743 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11540 18846 11552
rect 19245 11543 19303 11549
rect 19245 11540 19257 11543
rect 18840 11512 19257 11540
rect 18840 11500 18846 11512
rect 19245 11509 19257 11512
rect 19291 11540 19303 11543
rect 19518 11540 19524 11552
rect 19291 11512 19524 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 19610 11500 19616 11552
rect 19668 11540 19674 11552
rect 19886 11540 19892 11552
rect 19668 11512 19892 11540
rect 19668 11500 19674 11512
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 13814 11336 13820 11348
rect 11379 11308 13820 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 14608 11308 17325 11336
rect 14608 11296 14614 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 21174 11336 21180 11348
rect 21135 11308 21180 11336
rect 17313 11299 17371 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 14093 11271 14151 11277
rect 14093 11237 14105 11271
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 20717 11271 20775 11277
rect 20717 11237 20729 11271
rect 20763 11268 20775 11271
rect 20806 11268 20812 11280
rect 20763 11240 20812 11268
rect 20763 11237 20775 11240
rect 20717 11231 20775 11237
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 11698 11132 11704 11144
rect 9999 11104 11704 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 11698 11092 11704 11104
rect 11756 11132 11762 11144
rect 12342 11132 12348 11144
rect 11756 11104 12348 11132
rect 11756 11092 11762 11104
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 14108 11132 14136 11231
rect 20806 11228 20812 11240
rect 20864 11228 20870 11280
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 12492 11104 14136 11132
rect 15120 11104 15485 11132
rect 12492 11092 12498 11104
rect 10220 11067 10278 11073
rect 10220 11033 10232 11067
rect 10266 11064 10278 11067
rect 12544 11064 12572 11104
rect 15120 11076 15148 11104
rect 15473 11101 15485 11104
rect 15519 11132 15531 11135
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15519 11104 15761 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 18782 11132 18788 11144
rect 18739 11104 18788 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 18782 11092 18788 11104
rect 18840 11132 18846 11144
rect 19337 11135 19395 11141
rect 19337 11132 19349 11135
rect 18840 11104 19349 11132
rect 18840 11092 18846 11104
rect 19337 11101 19349 11104
rect 19383 11132 19395 11135
rect 21358 11132 21364 11144
rect 19383 11104 19840 11132
rect 21319 11104 21364 11132
rect 19383 11101 19395 11104
rect 19337 11095 19395 11101
rect 19812 11076 19840 11104
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 10266 11036 12572 11064
rect 12612 11067 12670 11073
rect 10266 11033 10278 11036
rect 10220 11027 10278 11033
rect 12612 11033 12624 11067
rect 12658 11064 12670 11067
rect 12986 11064 12992 11076
rect 12658 11036 12992 11064
rect 12658 11033 12670 11036
rect 12612 11027 12670 11033
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 15102 11024 15108 11076
rect 15160 11024 15166 11076
rect 15206 11067 15264 11073
rect 15206 11033 15218 11067
rect 15252 11033 15264 11067
rect 15206 11027 15264 11033
rect 13722 10996 13728 11008
rect 13683 10968 13728 10996
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 15010 10956 15016 11008
rect 15068 10996 15074 11008
rect 15212 10996 15240 11027
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18426 11067 18484 11073
rect 18426 11064 18438 11067
rect 18380 11036 18438 11064
rect 18380 11024 18386 11036
rect 18426 11033 18438 11036
rect 18472 11033 18484 11067
rect 18426 11027 18484 11033
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19582 11067 19640 11073
rect 19582 11064 19594 11067
rect 19116 11036 19594 11064
rect 19116 11024 19122 11036
rect 19582 11033 19594 11036
rect 19628 11033 19640 11067
rect 19582 11027 19640 11033
rect 19794 11024 19800 11076
rect 19852 11024 19858 11076
rect 15068 10968 15240 10996
rect 15068 10956 15074 10968
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 1636 10764 7389 10792
rect 1636 10752 1642 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 18230 10792 18236 10804
rect 7377 10755 7435 10761
rect 18064 10764 18236 10792
rect 12342 10724 12348 10736
rect 9692 10696 12348 10724
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 8018 10656 8024 10668
rect 7515 10628 8024 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 9692 10665 9720 10696
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 9944 10659 10002 10665
rect 9944 10656 9956 10659
rect 9824 10628 9956 10656
rect 9824 10616 9830 10628
rect 9944 10625 9956 10628
rect 9990 10656 10002 10659
rect 10870 10656 10876 10668
rect 9990 10628 10876 10656
rect 9990 10625 10002 10628
rect 9944 10619 10002 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11624 10665 11652 10696
rect 12342 10684 12348 10696
rect 12400 10724 12406 10736
rect 15102 10724 15108 10736
rect 12400 10684 12434 10724
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11865 10659 11923 10665
rect 11865 10656 11877 10659
rect 11609 10619 11667 10625
rect 11716 10628 11877 10656
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 8202 10588 8208 10600
rect 7331 10560 8208 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 11716 10588 11744 10628
rect 11865 10625 11877 10628
rect 11911 10625 11923 10659
rect 12406 10656 12434 10684
rect 13648 10696 15108 10724
rect 13648 10665 13676 10696
rect 15102 10684 15108 10696
rect 15160 10684 15166 10736
rect 16936 10727 16994 10733
rect 16936 10693 16948 10727
rect 16982 10724 16994 10727
rect 18064 10724 18092 10764
rect 18230 10752 18236 10764
rect 18288 10792 18294 10804
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 18288 10764 19993 10792
rect 18288 10752 18294 10764
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 16982 10696 18092 10724
rect 16982 10693 16994 10696
rect 16936 10687 16994 10693
rect 13357 10659 13415 10665
rect 13357 10656 13369 10659
rect 12406 10628 13369 10656
rect 11865 10619 11923 10625
rect 13357 10625 13369 10628
rect 13403 10656 13415 10659
rect 13633 10659 13691 10665
rect 13633 10656 13645 10659
rect 13403 10628 13645 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 13633 10625 13645 10628
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 13889 10659 13947 10665
rect 13889 10656 13901 10659
rect 13780 10628 13901 10656
rect 13780 10616 13786 10628
rect 13889 10625 13901 10628
rect 13935 10625 13947 10659
rect 19438 10659 19496 10665
rect 19438 10656 19450 10659
rect 13889 10619 13947 10625
rect 18064 10628 19450 10656
rect 11072 10560 11744 10588
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10520 7895 10523
rect 8294 10520 8300 10532
rect 7883 10492 8300 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 8076 10424 8125 10452
rect 8076 10412 8082 10424
rect 8113 10421 8125 10424
rect 8159 10421 8171 10455
rect 8113 10415 8171 10421
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 11072 10461 11100 10560
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 13740 10588 13768 10616
rect 12952 10560 13768 10588
rect 12952 10548 12958 10560
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 15160 10560 15393 10588
rect 15160 10548 15166 10560
rect 15381 10557 15393 10560
rect 15427 10588 15439 10591
rect 16666 10588 16672 10600
rect 15427 10560 16672 10588
rect 15427 10557 15439 10560
rect 15381 10551 15439 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 17862 10480 17868 10532
rect 17920 10520 17926 10532
rect 18064 10529 18092 10628
rect 19438 10625 19450 10628
rect 19484 10625 19496 10659
rect 19438 10619 19496 10625
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 19794 10656 19800 10668
rect 19751 10628 19800 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 19794 10616 19800 10628
rect 19852 10616 19858 10668
rect 20916 10656 20944 10752
rect 21266 10684 21272 10736
rect 21324 10724 21330 10736
rect 21324 10696 21404 10724
rect 21324 10684 21330 10696
rect 21376 10665 21404 10696
rect 21105 10659 21163 10665
rect 21105 10656 21117 10659
rect 20916 10628 21117 10656
rect 21105 10625 21117 10628
rect 21151 10656 21163 10659
rect 21361 10659 21419 10665
rect 21151 10628 21312 10656
rect 21151 10625 21163 10628
rect 21105 10619 21163 10625
rect 21284 10588 21312 10628
rect 21361 10625 21373 10659
rect 21407 10625 21419 10659
rect 21361 10619 21419 10625
rect 21542 10588 21548 10600
rect 21284 10560 21548 10588
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 17920 10492 18061 10520
rect 17920 10480 17926 10492
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 11020 10424 11069 10452
rect 11020 10412 11026 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 11057 10415 11115 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 15010 10452 15016 10464
rect 14424 10424 15016 10452
rect 14424 10412 14430 10424
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 9692 10220 11437 10248
rect 9692 10121 9720 10220
rect 11425 10217 11437 10220
rect 11471 10248 11483 10251
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11471 10220 11805 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 11793 10217 11805 10220
rect 11839 10248 11851 10251
rect 12342 10248 12348 10260
rect 11839 10220 12348 10248
rect 11839 10217 11851 10220
rect 11793 10211 11851 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 15102 10248 15108 10260
rect 14752 10220 15108 10248
rect 11057 10183 11115 10189
rect 11057 10149 11069 10183
rect 11103 10180 11115 10183
rect 11882 10180 11888 10192
rect 11103 10152 11888 10180
rect 11103 10149 11115 10152
rect 11057 10143 11115 10149
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 14752 10121 14780 10220
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 20070 10248 20076 10260
rect 20031 10220 20076 10248
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20809 10183 20867 10189
rect 20809 10180 20821 10183
rect 17696 10152 20821 10180
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 17696 10044 17724 10152
rect 20809 10149 20821 10152
rect 20855 10149 20867 10183
rect 20809 10143 20867 10149
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19576 10084 21036 10112
rect 19576 10072 19582 10084
rect 14516 10016 17724 10044
rect 18877 10047 18935 10053
rect 14516 10004 14522 10016
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19886 10044 19892 10056
rect 18923 10016 19892 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 20346 10044 20352 10056
rect 20307 10016 20352 10044
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 21008 10053 21036 10084
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 9950 9985 9956 9988
rect 9944 9939 9956 9985
rect 10008 9976 10014 9988
rect 10008 9948 10044 9976
rect 9950 9936 9956 9939
rect 10008 9936 10014 9948
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 14982 9979 15040 9985
rect 14982 9976 14994 9979
rect 13872 9948 14994 9976
rect 13872 9936 13878 9948
rect 14982 9945 14994 9948
rect 15028 9945 15040 9979
rect 14982 9939 15040 9945
rect 16485 9979 16543 9985
rect 16485 9945 16497 9979
rect 16531 9976 16543 9979
rect 16666 9976 16672 9988
rect 16531 9948 16672 9976
rect 16531 9945 16543 9948
rect 16485 9939 16543 9945
rect 16666 9936 16672 9948
rect 16724 9976 16730 9988
rect 18233 9979 18291 9985
rect 18233 9976 18245 9979
rect 16724 9948 18245 9976
rect 16724 9936 16730 9948
rect 18233 9945 18245 9948
rect 18279 9976 18291 9979
rect 19613 9979 19671 9985
rect 19613 9976 19625 9979
rect 18279 9948 19625 9976
rect 18279 9945 18291 9948
rect 18233 9939 18291 9945
rect 19613 9945 19625 9948
rect 19659 9976 19671 9979
rect 19794 9976 19800 9988
rect 19659 9948 19800 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 19794 9936 19800 9948
rect 19852 9976 19858 9988
rect 19852 9948 21312 9976
rect 19852 9936 19858 9948
rect 21284 9920 21312 9948
rect 20530 9908 20536 9920
rect 20491 9880 20536 9908
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 21266 9908 21272 9920
rect 21227 9880 21272 9908
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 8205 9707 8263 9713
rect 8205 9673 8217 9707
rect 8251 9704 8263 9707
rect 8294 9704 8300 9716
rect 8251 9676 8300 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 19061 9707 19119 9713
rect 19061 9673 19073 9707
rect 19107 9704 19119 9707
rect 20346 9704 20352 9716
rect 19107 9676 20352 9704
rect 19107 9673 19119 9676
rect 19061 9667 19119 9673
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 10410 9596 10416 9648
rect 10468 9636 10474 9648
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 10468 9608 11529 9636
rect 10468 9596 10474 9608
rect 11517 9605 11529 9608
rect 11563 9636 11575 9639
rect 18138 9636 18144 9648
rect 11563 9608 18144 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 18325 9639 18383 9645
rect 18325 9605 18337 9639
rect 18371 9636 18383 9639
rect 18414 9636 18420 9648
rect 18371 9608 18420 9636
rect 18371 9605 18383 9608
rect 18325 9599 18383 9605
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 18693 9639 18751 9645
rect 18693 9605 18705 9639
rect 18739 9636 18751 9639
rect 18739 9608 20944 9636
rect 18739 9605 18751 9608
rect 18693 9599 18751 9605
rect 20916 9580 20944 9608
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8570 9568 8576 9580
rect 8343 9540 8576 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 9398 9528 9404 9580
rect 9456 9568 9462 9580
rect 13538 9568 13544 9580
rect 9456 9540 13544 9568
rect 9456 9528 9462 9540
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 19337 9571 19395 9577
rect 19337 9537 19349 9571
rect 19383 9568 19395 9571
rect 19794 9568 19800 9580
rect 19383 9540 19800 9568
rect 19383 9537 19395 9540
rect 19337 9531 19395 9537
rect 19794 9528 19800 9540
rect 19852 9528 19858 9580
rect 19981 9571 20039 9577
rect 19981 9537 19993 9571
rect 20027 9537 20039 9571
rect 20254 9568 20260 9580
rect 20215 9540 20260 9568
rect 19981 9531 20039 9537
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 10870 9500 10876 9512
rect 8159 9472 10876 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 19996 9500 20024 9531
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20898 9568 20904 9580
rect 20859 9540 20904 9568
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 21174 9568 21180 9580
rect 21135 9540 21180 9568
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 20990 9500 20996 9512
rect 19996 9472 20996 9500
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 14642 9432 14648 9444
rect 7892 9404 14648 9432
rect 7892 9392 7898 9404
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 19521 9435 19579 9441
rect 19521 9401 19533 9435
rect 19567 9432 19579 9435
rect 19978 9432 19984 9444
rect 19567 9404 19984 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 19978 9392 19984 9404
rect 20036 9392 20042 9444
rect 20438 9432 20444 9444
rect 20399 9404 20444 9432
rect 20438 9392 20444 9404
rect 20496 9392 20502 9444
rect 20714 9432 20720 9444
rect 20675 9404 20720 9432
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 21361 9435 21419 9441
rect 21361 9401 21373 9435
rect 21407 9432 21419 9435
rect 21450 9432 21456 9444
rect 21407 9404 21456 9432
rect 21407 9401 21419 9404
rect 21361 9395 21419 9401
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 10686 9364 10692 9376
rect 8711 9336 10692 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 15378 9364 15384 9376
rect 15339 9336 15384 9364
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 16264 9336 19809 9364
rect 16264 9324 16270 9336
rect 19797 9333 19809 9336
rect 19843 9333 19855 9367
rect 19797 9327 19855 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 8570 9160 8576 9172
rect 8531 9132 8576 9160
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 10560 9132 11437 9160
rect 10560 9120 10566 9132
rect 11425 9129 11437 9132
rect 11471 9129 11483 9163
rect 17681 9163 17739 9169
rect 17681 9160 17693 9163
rect 11425 9123 11483 9129
rect 11716 9132 17693 9160
rect 10962 9092 10968 9104
rect 10520 9064 10968 9092
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8202 9024 8208 9036
rect 8067 8996 8208 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 10520 9033 10548 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10686 9024 10692 9036
rect 10647 8996 10692 9024
rect 10505 8987 10563 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 11716 8956 11744 9132
rect 17681 9129 17693 9132
rect 17727 9129 17739 9163
rect 17681 9123 17739 9129
rect 19429 9163 19487 9169
rect 19429 9129 19441 9163
rect 19475 9160 19487 9163
rect 20254 9160 20260 9172
rect 19475 9132 20260 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 21082 9160 21088 9172
rect 21043 9132 21088 9160
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 11882 9052 11888 9104
rect 11940 9092 11946 9104
rect 13449 9095 13507 9101
rect 11940 9064 12020 9092
rect 11940 9052 11946 9064
rect 11992 9033 12020 9064
rect 13449 9061 13461 9095
rect 13495 9092 13507 9095
rect 17405 9095 17463 9101
rect 13495 9064 15792 9092
rect 13495 9061 13507 9064
rect 13449 9055 13507 9061
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 9024 12955 9027
rect 13814 9024 13820 9036
rect 12943 8996 13820 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 13814 8984 13820 8996
rect 13872 9024 13878 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 13872 8996 14565 9024
rect 13872 8984 13878 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14553 8987 14611 8993
rect 14660 8996 14749 9024
rect 8168 8928 11744 8956
rect 8168 8916 8174 8928
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 8128 8860 8953 8888
rect 7834 8780 7840 8832
rect 7892 8820 7898 8832
rect 8128 8829 8156 8860
rect 8941 8857 8953 8860
rect 8987 8857 8999 8891
rect 8941 8851 8999 8857
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 11885 8891 11943 8897
rect 11885 8888 11897 8891
rect 10468 8860 11897 8888
rect 10468 8848 10474 8860
rect 11885 8857 11897 8860
rect 11931 8857 11943 8891
rect 11885 8851 11943 8857
rect 12066 8848 12072 8900
rect 12124 8888 12130 8900
rect 14660 8888 14688 8996
rect 14737 8993 14749 8996
rect 14783 9024 14795 9027
rect 15378 9024 15384 9036
rect 14783 8996 15384 9024
rect 14783 8993 14795 8996
rect 14737 8987 14795 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15764 9033 15792 9064
rect 17405 9061 17417 9095
rect 17451 9092 17463 9095
rect 17451 9064 21312 9092
rect 17451 9061 17463 9064
rect 17405 9055 17463 9061
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 19058 9024 19064 9036
rect 18371 8996 19064 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 15672 8956 15700 8987
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 19794 9024 19800 9036
rect 19755 8996 19800 9024
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 20622 9024 20628 9036
rect 20583 8996 20628 9024
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 16114 8956 16120 8968
rect 15672 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 17221 8959 17279 8965
rect 17221 8956 17233 8959
rect 17184 8928 17233 8956
rect 17184 8916 17190 8928
rect 17221 8925 17233 8928
rect 17267 8925 17279 8959
rect 19242 8956 19248 8968
rect 17221 8919 17279 8925
rect 17328 8928 18828 8956
rect 19203 8928 19248 8956
rect 15841 8891 15899 8897
rect 15841 8888 15853 8891
rect 12124 8860 14688 8888
rect 15212 8860 15853 8888
rect 12124 8848 12130 8860
rect 8113 8823 8171 8829
rect 8113 8820 8125 8823
rect 7892 8792 8125 8820
rect 7892 8780 7898 8792
rect 8113 8789 8125 8792
rect 8159 8789 8171 8823
rect 8113 8783 8171 8789
rect 8205 8823 8263 8829
rect 8205 8789 8217 8823
rect 8251 8820 8263 8823
rect 9398 8820 9404 8832
rect 8251 8792 9404 8820
rect 8251 8789 8263 8792
rect 8205 8783 8263 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11146 8820 11152 8832
rect 10836 8792 10881 8820
rect 11107 8792 11152 8820
rect 10836 8780 10842 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11790 8820 11796 8832
rect 11751 8792 11796 8820
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12308 8792 13001 8820
rect 12308 8780 12314 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 12989 8783 13047 8789
rect 13081 8823 13139 8829
rect 13081 8789 13093 8823
rect 13127 8820 13139 8823
rect 13170 8820 13176 8832
rect 13127 8792 13176 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 14185 8823 14243 8829
rect 14185 8820 14197 8823
rect 13596 8792 14197 8820
rect 13596 8780 13602 8792
rect 14185 8789 14197 8792
rect 14231 8820 14243 8823
rect 14458 8820 14464 8832
rect 14231 8792 14464 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14829 8823 14887 8829
rect 14829 8789 14841 8823
rect 14875 8820 14887 8823
rect 14918 8820 14924 8832
rect 14875 8792 14924 8820
rect 14875 8789 14887 8792
rect 14829 8783 14887 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 15212 8829 15240 8860
rect 15841 8857 15853 8860
rect 15887 8857 15899 8891
rect 15841 8851 15899 8857
rect 16298 8848 16304 8900
rect 16356 8888 16362 8900
rect 17328 8888 17356 8928
rect 16356 8860 17356 8888
rect 18049 8891 18107 8897
rect 16356 8848 16362 8860
rect 18049 8857 18061 8891
rect 18095 8888 18107 8891
rect 18693 8891 18751 8897
rect 18693 8888 18705 8891
rect 18095 8860 18705 8888
rect 18095 8857 18107 8860
rect 18049 8851 18107 8857
rect 18693 8857 18705 8860
rect 18739 8857 18751 8891
rect 18800 8888 18828 8928
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 20441 8959 20499 8965
rect 20441 8925 20453 8959
rect 20487 8956 20499 8959
rect 20530 8956 20536 8968
rect 20487 8928 20536 8956
rect 20487 8925 20499 8928
rect 20441 8919 20499 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 21284 8965 21312 9064
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 22094 8888 22100 8900
rect 18800 8860 22100 8888
rect 18693 8851 18751 8857
rect 22094 8848 22100 8860
rect 22152 8848 22158 8900
rect 15197 8823 15255 8829
rect 15197 8789 15209 8823
rect 15243 8789 15255 8823
rect 16206 8820 16212 8832
rect 16167 8792 16212 8820
rect 15197 8783 15255 8789
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 19058 8820 19064 8832
rect 18187 8792 19064 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 20070 8820 20076 8832
rect 20031 8792 20076 8820
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 20530 8820 20536 8832
rect 20491 8792 20536 8820
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10778 8616 10784 8628
rect 10459 8588 10784 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 12250 8616 12256 8628
rect 11204 8588 12112 8616
rect 12211 8588 12256 8616
rect 11204 8576 11210 8588
rect 11698 8548 11704 8560
rect 6886 8520 11704 8548
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 6886 8412 6914 8520
rect 11698 8508 11704 8520
rect 11756 8548 11762 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11756 8520 11805 8548
rect 11756 8508 11762 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 12084 8548 12112 8588
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13538 8616 13544 8628
rect 13499 8588 13544 8616
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13633 8619 13691 8625
rect 13633 8585 13645 8619
rect 13679 8616 13691 8619
rect 14642 8616 14648 8628
rect 13679 8588 14648 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 14918 8616 14924 8628
rect 14879 8588 14924 8616
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 16298 8616 16304 8628
rect 16255 8588 16304 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 16669 8619 16727 8625
rect 16669 8585 16681 8619
rect 16715 8585 16727 8619
rect 17126 8616 17132 8628
rect 17087 8588 17132 8616
rect 16669 8579 16727 8585
rect 12084 8520 14228 8548
rect 11793 8511 11851 8517
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11238 8480 11244 8492
rect 10827 8452 11244 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 14200 8489 14228 8520
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 15286 8548 15292 8560
rect 14516 8520 15292 8548
rect 14516 8508 14522 8520
rect 15286 8508 15292 8520
rect 15344 8508 15350 8560
rect 16684 8548 16712 8579
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18196 8588 18705 8616
rect 18196 8576 18202 8588
rect 18693 8585 18705 8588
rect 18739 8616 18751 8619
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 18739 8588 19533 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 19521 8585 19533 8588
rect 19567 8616 19579 8619
rect 19886 8616 19892 8628
rect 19567 8588 19892 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 19886 8576 19892 8588
rect 19944 8616 19950 8628
rect 20530 8616 20536 8628
rect 19944 8588 20536 8616
rect 19944 8576 19950 8588
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 20809 8619 20867 8625
rect 20809 8585 20821 8619
rect 20855 8585 20867 8619
rect 21266 8616 21272 8628
rect 21227 8588 21272 8616
rect 20809 8579 20867 8585
rect 20824 8548 20852 8579
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 16040 8520 16712 8548
rect 17328 8520 20852 8548
rect 16040 8489 16068 8520
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11348 8452 11897 8480
rect 2372 8384 6914 8412
rect 2372 8372 2378 8384
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 10870 8412 10876 8424
rect 10744 8384 10876 8412
rect 10744 8372 10750 8384
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11020 8384 11065 8412
rect 11020 8372 11026 8384
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 11348 8344 11376 8452
rect 11885 8449 11897 8452
rect 11931 8480 11943 8483
rect 14185 8483 14243 8489
rect 11931 8452 12664 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 12434 8412 12440 8424
rect 11747 8384 12440 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12636 8421 12664 8452
rect 13648 8452 14136 8480
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8412 12679 8415
rect 13648 8412 13676 8452
rect 12667 8384 13676 8412
rect 13725 8415 13783 8421
rect 12667 8381 12679 8384
rect 12621 8375 12679 8381
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 14108 8412 14136 8452
rect 14185 8449 14197 8483
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16264 8452 16865 8480
rect 16264 8440 16270 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 14108 8384 15424 8412
rect 13725 8375 13783 8381
rect 8076 8316 11376 8344
rect 12452 8344 12480 8372
rect 13740 8344 13768 8375
rect 12452 8316 13768 8344
rect 14369 8347 14427 8353
rect 8076 8304 8082 8316
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 15194 8344 15200 8356
rect 14415 8316 15200 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 15396 8344 15424 8384
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 17328 8412 17356 8520
rect 17494 8480 17500 8492
rect 17455 8452 17500 8480
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 19794 8480 19800 8492
rect 19475 8452 19800 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20346 8480 20352 8492
rect 20307 8452 20352 8480
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20990 8480 20996 8492
rect 20951 8452 20996 8480
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 15528 8384 17356 8412
rect 15528 8372 15534 8384
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 17460 8384 17601 8412
rect 17460 8372 17466 8384
rect 17589 8381 17601 8384
rect 17635 8381 17647 8415
rect 17589 8375 17647 8381
rect 17773 8415 17831 8421
rect 17773 8381 17785 8415
rect 17819 8412 17831 8415
rect 18322 8412 18328 8424
rect 17819 8384 18328 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 19613 8415 19671 8421
rect 19613 8381 19625 8415
rect 19659 8381 19671 8415
rect 19613 8375 19671 8381
rect 17954 8344 17960 8356
rect 15396 8316 17960 8344
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 19628 8344 19656 8375
rect 18932 8316 19656 8344
rect 20533 8347 20591 8353
rect 18932 8304 18938 8316
rect 20533 8313 20545 8347
rect 20579 8344 20591 8347
rect 20898 8344 20904 8356
rect 20579 8316 20904 8344
rect 20579 8313 20591 8316
rect 20533 8307 20591 8313
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 19058 8276 19064 8288
rect 19019 8248 19064 8276
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 21634 8276 21640 8288
rect 20772 8248 21640 8276
rect 20772 8236 20778 8248
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 17405 8075 17463 8081
rect 17405 8041 17417 8075
rect 17451 8072 17463 8075
rect 17494 8072 17500 8084
rect 17451 8044 17500 8072
rect 17451 8041 17463 8044
rect 17405 8035 17463 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 20346 8072 20352 8084
rect 19659 8044 20352 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 20441 8075 20499 8081
rect 20441 8041 20453 8075
rect 20487 8072 20499 8075
rect 20990 8072 20996 8084
rect 20487 8044 20996 8072
rect 20487 8041 20499 8044
rect 20441 8035 20499 8041
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 12066 8004 12072 8016
rect 11112 7976 12072 8004
rect 11112 7964 11118 7976
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 14277 8007 14335 8013
rect 14277 7973 14289 8007
rect 14323 7973 14335 8007
rect 14277 7967 14335 7973
rect 15565 8007 15623 8013
rect 15565 7973 15577 8007
rect 15611 8004 15623 8007
rect 20530 8004 20536 8016
rect 15611 7976 20536 8004
rect 15611 7973 15623 7976
rect 15565 7967 15623 7973
rect 11238 7936 11244 7948
rect 11199 7908 11244 7936
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 14292 7936 14320 7967
rect 20530 7964 20536 7976
rect 20588 7964 20594 8016
rect 20714 8004 20720 8016
rect 20675 7976 20720 8004
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 22278 8004 22284 8016
rect 21232 7976 22284 8004
rect 21232 7964 21238 7976
rect 22278 7964 22284 7976
rect 22336 7964 22342 8016
rect 14292 7908 17816 7936
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13872 7840 14105 7868
rect 13872 7828 13878 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15252 7840 15393 7868
rect 15252 7828 15258 7840
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 17788 7868 17816 7908
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 17957 7939 18015 7945
rect 17957 7936 17969 7939
rect 17920 7908 17969 7936
rect 17920 7896 17926 7908
rect 17957 7905 17969 7908
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 19242 7896 19248 7948
rect 19300 7936 19306 7948
rect 19300 7908 21404 7936
rect 19300 7896 19306 7908
rect 21376 7880 21404 7908
rect 20257 7871 20315 7877
rect 17788 7840 18552 7868
rect 15381 7831 15439 7837
rect 17773 7803 17831 7809
rect 17773 7769 17785 7803
rect 17819 7800 17831 7803
rect 18417 7803 18475 7809
rect 18417 7800 18429 7803
rect 17819 7772 18429 7800
rect 17819 7769 17831 7772
rect 17773 7763 17831 7769
rect 18417 7769 18429 7772
rect 18463 7769 18475 7803
rect 18417 7763 18475 7769
rect 14642 7732 14648 7744
rect 14555 7704 14648 7732
rect 14642 7692 14648 7704
rect 14700 7732 14706 7744
rect 15010 7732 15016 7744
rect 14700 7704 15016 7732
rect 14700 7692 14706 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 17862 7732 17868 7744
rect 17823 7704 17868 7732
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 18524 7732 18552 7840
rect 20257 7837 20269 7871
rect 20303 7837 20315 7871
rect 20898 7868 20904 7880
rect 20859 7840 20904 7868
rect 20257 7831 20315 7837
rect 19886 7800 19892 7812
rect 19847 7772 19892 7800
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 20272 7800 20300 7831
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21174 7868 21180 7880
rect 21048 7840 21180 7868
rect 21048 7828 21054 7840
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21358 7868 21364 7880
rect 21319 7840 21364 7868
rect 21358 7828 21364 7840
rect 21416 7828 21422 7880
rect 20272 7772 21404 7800
rect 21376 7744 21404 7772
rect 20990 7732 20996 7744
rect 18524 7704 20996 7732
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 21174 7732 21180 7744
rect 21135 7704 21180 7732
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 21358 7692 21364 7744
rect 21416 7692 21422 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 19242 7528 19248 7540
rect 19203 7500 19248 7528
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7528 20039 7531
rect 20070 7528 20076 7540
rect 20027 7500 20076 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 21140 7500 21189 7528
rect 21140 7488 21146 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 11977 7463 12035 7469
rect 11977 7460 11989 7463
rect 11940 7432 11989 7460
rect 11940 7420 11946 7432
rect 11977 7429 11989 7432
rect 12023 7429 12035 7463
rect 11977 7423 12035 7429
rect 18877 7463 18935 7469
rect 18877 7429 18889 7463
rect 18923 7460 18935 7463
rect 18923 7432 21404 7460
rect 18923 7429 18935 7432
rect 18877 7423 18935 7429
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 21376 7401 21404 7432
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 2924 7364 11069 7392
rect 2924 7352 2930 7364
rect 11057 7361 11069 7364
rect 11103 7392 11115 7395
rect 19889 7395 19947 7401
rect 11103 7364 11928 7392
rect 11103 7361 11115 7364
rect 11057 7355 11115 7361
rect 11900 7333 11928 7364
rect 19889 7361 19901 7395
rect 19935 7392 19947 7395
rect 20533 7395 20591 7401
rect 20533 7392 20545 7395
rect 19935 7364 20545 7392
rect 19935 7361 19947 7364
rect 19889 7355 19947 7361
rect 20533 7361 20545 7364
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21450 7392 21456 7404
rect 21407 7364 21456 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 11793 7327 11851 7333
rect 11793 7293 11805 7327
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 11885 7327 11943 7333
rect 11885 7293 11897 7327
rect 11931 7293 11943 7327
rect 11885 7287 11943 7293
rect 20073 7327 20131 7333
rect 20073 7293 20085 7327
rect 20119 7324 20131 7327
rect 21542 7324 21548 7336
rect 20119 7296 21548 7324
rect 20119 7293 20131 7296
rect 20073 7287 20131 7293
rect 11808 7256 11836 7287
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 14274 7256 14280 7268
rect 11808 7228 14280 7256
rect 14274 7216 14280 7228
rect 14332 7256 14338 7268
rect 14918 7256 14924 7268
rect 14332 7228 14924 7256
rect 14332 7216 14338 7228
rect 14918 7216 14924 7228
rect 14976 7216 14982 7268
rect 19521 7259 19579 7265
rect 19521 7225 19533 7259
rect 19567 7256 19579 7259
rect 20162 7256 20168 7268
rect 19567 7228 20168 7256
rect 19567 7225 19579 7228
rect 19521 7219 19579 7225
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 12345 7191 12403 7197
rect 12345 7157 12357 7191
rect 12391 7188 12403 7191
rect 13630 7188 13636 7200
rect 12391 7160 13636 7188
rect 12391 7157 12403 7160
rect 12345 7151 12403 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 15194 7188 15200 7200
rect 15107 7160 15200 7188
rect 15194 7148 15200 7160
rect 15252 7188 15258 7200
rect 15930 7188 15936 7200
rect 15252 7160 15936 7188
rect 15252 7148 15258 7160
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 13688 6820 14596 6848
rect 13688 6808 13694 6820
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13722 6780 13728 6792
rect 13495 6752 13728 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 14568 6780 14596 6820
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 14700 6820 14745 6848
rect 14700 6808 14706 6820
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 15473 6851 15531 6857
rect 15473 6848 15485 6851
rect 14976 6820 15485 6848
rect 14976 6808 14982 6820
rect 15473 6817 15485 6820
rect 15519 6817 15531 6851
rect 15473 6811 15531 6817
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 17034 6848 17040 6860
rect 16623 6820 17040 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17828 6820 17969 6848
rect 17828 6808 17834 6820
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 19610 6808 19616 6860
rect 19668 6848 19674 6860
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19668 6820 19809 6848
rect 19668 6808 19674 6820
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 19797 6811 19855 6817
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 21358 6848 21364 6860
rect 20036 6820 21036 6848
rect 21319 6820 21364 6848
rect 20036 6808 20042 6820
rect 16669 6783 16727 6789
rect 16669 6780 16681 6783
rect 14568 6752 16681 6780
rect 16669 6749 16681 6752
rect 16715 6749 16727 6783
rect 20346 6780 20352 6792
rect 20307 6752 20352 6780
rect 16669 6743 16727 6749
rect 20346 6740 20352 6752
rect 20404 6740 20410 6792
rect 21008 6789 21036 6820
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 14553 6715 14611 6721
rect 9180 6684 14504 6712
rect 9180 6672 9186 6684
rect 13633 6647 13691 6653
rect 13633 6613 13645 6647
rect 13679 6644 13691 6647
rect 13814 6644 13820 6656
rect 13679 6616 13820 6644
rect 13679 6613 13691 6616
rect 13633 6607 13691 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 14476 6653 14504 6684
rect 14553 6681 14565 6715
rect 14599 6712 14611 6715
rect 14826 6712 14832 6724
rect 14599 6684 14832 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 16761 6715 16819 6721
rect 16761 6712 16773 6715
rect 16132 6684 16773 6712
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13964 6616 14105 6644
rect 13964 6604 13970 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 14461 6647 14519 6653
rect 14461 6613 14473 6647
rect 14507 6644 14519 6647
rect 15194 6644 15200 6656
rect 14507 6616 15200 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15654 6644 15660 6656
rect 15615 6616 15660 6644
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 16132 6653 16160 6684
rect 16761 6681 16773 6684
rect 16807 6681 16819 6715
rect 16761 6675 16819 6681
rect 17494 6672 17500 6724
rect 17552 6712 17558 6724
rect 17865 6715 17923 6721
rect 17865 6712 17877 6715
rect 17552 6684 17877 6712
rect 17552 6672 17558 6684
rect 17865 6681 17877 6684
rect 17911 6681 17923 6715
rect 17865 6675 17923 6681
rect 18877 6715 18935 6721
rect 18877 6681 18889 6715
rect 18923 6712 18935 6715
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 18923 6684 19625 6712
rect 18923 6681 18935 6684
rect 18877 6675 18935 6681
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 16117 6647 16175 6653
rect 15804 6616 15849 6644
rect 15804 6604 15810 6616
rect 16117 6613 16129 6647
rect 16163 6613 16175 6647
rect 16117 6607 16175 6613
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17218 6644 17224 6656
rect 17175 6616 17224 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17678 6604 17684 6656
rect 17736 6644 17742 6656
rect 17773 6647 17831 6653
rect 17773 6644 17785 6647
rect 17736 6616 17785 6644
rect 17736 6604 17742 6616
rect 17773 6613 17785 6616
rect 17819 6613 17831 6647
rect 17773 6607 17831 6613
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 18104 6616 19257 6644
rect 18104 6604 18110 6616
rect 19245 6613 19257 6616
rect 19291 6613 19303 6647
rect 19245 6607 19303 6613
rect 19705 6647 19763 6653
rect 19705 6613 19717 6647
rect 19751 6644 19763 6647
rect 20254 6644 20260 6656
rect 19751 6616 20260 6644
rect 19751 6613 19763 6616
rect 19705 6607 19763 6613
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20533 6647 20591 6653
rect 20533 6613 20545 6647
rect 20579 6644 20591 6647
rect 20622 6644 20628 6656
rect 20579 6616 20628 6644
rect 20579 6613 20591 6616
rect 20533 6607 20591 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 20772 6616 20821 6644
rect 20772 6604 20778 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12989 6443 13047 6449
rect 12989 6440 13001 6443
rect 12299 6412 13001 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12989 6409 13001 6412
rect 13035 6409 13047 6443
rect 12989 6403 13047 6409
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13495 6412 14197 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 14921 6443 14979 6449
rect 14921 6440 14933 6443
rect 14884 6412 14933 6440
rect 14884 6400 14890 6412
rect 14921 6409 14933 6412
rect 14967 6409 14979 6443
rect 15746 6440 15752 6452
rect 15707 6412 15752 6440
rect 14921 6403 14979 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 17405 6443 17463 6449
rect 15988 6412 17264 6440
rect 15988 6400 15994 6412
rect 1762 6332 1768 6384
rect 1820 6372 1826 6384
rect 11057 6375 11115 6381
rect 11057 6372 11069 6375
rect 1820 6344 11069 6372
rect 1820 6332 1826 6344
rect 11057 6341 11069 6344
rect 11103 6372 11115 6375
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11103 6344 11805 6372
rect 11103 6341 11115 6344
rect 11057 6335 11115 6341
rect 11793 6341 11805 6344
rect 11839 6341 11851 6375
rect 11793 6335 11851 6341
rect 13081 6375 13139 6381
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13906 6372 13912 6384
rect 13127 6344 13912 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 15194 6372 15200 6384
rect 14016 6344 15200 6372
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6304 1458 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1452 6276 1869 6304
rect 1452 6264 1458 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 11882 6304 11888 6316
rect 11795 6276 11888 6304
rect 1857 6267 1915 6273
rect 11882 6264 11888 6276
rect 11940 6304 11946 6316
rect 14016 6304 14044 6344
rect 15194 6332 15200 6344
rect 15252 6372 15258 6384
rect 17037 6375 17095 6381
rect 17037 6372 17049 6375
rect 15252 6344 17049 6372
rect 15252 6332 15258 6344
rect 17037 6341 17049 6344
rect 17083 6341 17095 6375
rect 17037 6335 17095 6341
rect 11940 6276 14044 6304
rect 14093 6307 14151 6313
rect 11940 6264 11946 6276
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 15102 6304 15108 6316
rect 14139 6276 15108 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 17236 6304 17264 6412
rect 17405 6409 17417 6443
rect 17451 6440 17463 6443
rect 17494 6440 17500 6452
rect 17451 6412 17500 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 17678 6440 17684 6452
rect 17639 6412 17684 6440
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 19518 6440 19524 6452
rect 19479 6412 19524 6440
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 20254 6440 20260 6452
rect 20215 6412 20260 6440
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 20622 6440 20628 6452
rect 20583 6412 20628 6440
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 21358 6440 21364 6452
rect 21319 6412 21364 6440
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 17310 6332 17316 6384
rect 17368 6372 17374 6384
rect 17368 6344 19840 6372
rect 17368 6332 17374 6344
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 16868 6276 17071 6304
rect 17236 6276 18061 6304
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6205 11759 6239
rect 12894 6236 12900 6248
rect 12855 6208 12900 6236
rect 11701 6199 11759 6205
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 9950 6168 9956 6180
rect 1627 6140 9956 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 11716 6168 11744 6199
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 14366 6236 14372 6248
rect 13556 6208 13860 6236
rect 14327 6208 14372 6236
rect 12986 6168 12992 6180
rect 11716 6140 12992 6168
rect 12986 6128 12992 6140
rect 13044 6168 13050 6180
rect 13556 6168 13584 6208
rect 13722 6168 13728 6180
rect 13044 6140 13584 6168
rect 13683 6140 13728 6168
rect 13044 6128 13050 6140
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 13832 6168 13860 6208
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 16868 6245 16896 6276
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6205 17003 6239
rect 16945 6199 17003 6205
rect 14642 6168 14648 6180
rect 13832 6140 14648 6168
rect 14642 6128 14648 6140
rect 14700 6128 14706 6180
rect 16209 6171 16267 6177
rect 16209 6168 16221 6171
rect 14844 6140 16221 6168
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 14844 6100 14872 6140
rect 16209 6137 16221 6140
rect 16255 6168 16267 6171
rect 16960 6168 16988 6199
rect 16255 6140 16988 6168
rect 17043 6168 17071 6276
rect 18049 6273 18061 6276
rect 18095 6304 18107 6307
rect 18874 6304 18880 6316
rect 18095 6276 18460 6304
rect 18835 6276 18880 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 18138 6236 18144 6248
rect 18099 6208 18144 6236
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18230 6196 18236 6248
rect 18288 6236 18294 6248
rect 18288 6208 18333 6236
rect 18288 6196 18294 6208
rect 18248 6168 18276 6196
rect 17043 6140 18276 6168
rect 18432 6168 18460 6276
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19812 6313 19840 6344
rect 19886 6332 19892 6384
rect 19944 6372 19950 6384
rect 20530 6372 20536 6384
rect 19944 6344 20536 6372
rect 19944 6332 19950 6344
rect 20530 6332 20536 6344
rect 20588 6372 20594 6384
rect 20717 6375 20775 6381
rect 20717 6372 20729 6375
rect 20588 6344 20729 6372
rect 20588 6332 20594 6344
rect 20717 6341 20729 6344
rect 20763 6341 20775 6375
rect 20717 6335 20775 6341
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6273 19855 6307
rect 21376 6304 21404 6400
rect 19797 6267 19855 6273
rect 19904 6276 21404 6304
rect 19352 6236 19380 6267
rect 19904 6236 19932 6276
rect 19352 6208 19932 6236
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 20864 6208 20909 6236
rect 20864 6196 20870 6208
rect 19518 6168 19524 6180
rect 18432 6140 19524 6168
rect 16255 6137 16267 6140
rect 16209 6131 16267 6137
rect 19518 6128 19524 6140
rect 19576 6128 19582 6180
rect 12400 6072 14872 6100
rect 12400 6060 12406 6072
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 18138 6100 18144 6112
rect 14976 6072 18144 6100
rect 14976 6060 14982 6072
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 19058 6100 19064 6112
rect 19019 6072 19064 6100
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 19981 6103 20039 6109
rect 19981 6069 19993 6103
rect 20027 6100 20039 6103
rect 20806 6100 20812 6112
rect 20027 6072 20812 6100
rect 20027 6069 20039 6072
rect 19981 6063 20039 6069
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 17862 5896 17868 5908
rect 17819 5868 17868 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18782 5896 18788 5908
rect 18196 5868 18788 5896
rect 18196 5856 18202 5868
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 19794 5896 19800 5908
rect 19755 5868 19800 5896
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 20588 5868 21281 5896
rect 20588 5856 20594 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 17586 5788 17592 5840
rect 17644 5828 17650 5840
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 17644 5800 20269 5828
rect 17644 5788 17650 5800
rect 20257 5797 20269 5800
rect 20303 5797 20315 5831
rect 20714 5828 20720 5840
rect 20675 5800 20720 5828
rect 20257 5791 20315 5797
rect 20714 5788 20720 5800
rect 20772 5788 20778 5840
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 12952 5732 15669 5760
rect 12952 5720 12958 5732
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 18288 5732 18337 5760
rect 18288 5720 18294 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 19058 5720 19064 5772
rect 19116 5760 19122 5772
rect 19116 5732 20944 5760
rect 19116 5720 19122 5732
rect 19978 5692 19984 5704
rect 19939 5664 19984 5692
rect 19978 5652 19984 5664
rect 20036 5652 20042 5704
rect 20916 5701 20944 5732
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 15473 5627 15531 5633
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 16117 5627 16175 5633
rect 16117 5624 16129 5627
rect 15519 5596 16129 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 16117 5593 16129 5596
rect 16163 5593 16175 5627
rect 18322 5624 18328 5636
rect 16117 5587 16175 5593
rect 18156 5596 18328 5624
rect 15562 5556 15568 5568
rect 15523 5528 15568 5556
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 18156 5565 18184 5596
rect 18322 5584 18328 5596
rect 18380 5584 18386 5636
rect 20456 5624 20484 5655
rect 21174 5624 21180 5636
rect 20456 5596 21180 5624
rect 21174 5584 21180 5596
rect 21232 5584 21238 5636
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 19337 5559 19395 5565
rect 18288 5528 18333 5556
rect 18288 5516 18294 5528
rect 19337 5525 19349 5559
rect 19383 5556 19395 5559
rect 19518 5556 19524 5568
rect 19383 5528 19524 5556
rect 19383 5525 19395 5528
rect 19337 5519 19395 5525
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 15105 5355 15163 5361
rect 15105 5321 15117 5355
rect 15151 5352 15163 5355
rect 15562 5352 15568 5364
rect 15151 5324 15568 5352
rect 15151 5321 15163 5324
rect 15105 5315 15163 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 19242 5352 19248 5364
rect 19203 5324 19248 5352
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 19978 5352 19984 5364
rect 19659 5324 19984 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20346 5312 20352 5364
rect 20404 5352 20410 5364
rect 21269 5355 21327 5361
rect 21269 5352 21281 5355
rect 20404 5324 21281 5352
rect 20404 5312 20410 5324
rect 21269 5321 21281 5324
rect 21315 5321 21327 5355
rect 21269 5315 21327 5321
rect 15473 5287 15531 5293
rect 15473 5253 15485 5287
rect 15519 5284 15531 5287
rect 15654 5284 15660 5296
rect 15519 5256 15660 5284
rect 15519 5253 15531 5256
rect 15473 5247 15531 5253
rect 15654 5244 15660 5256
rect 15712 5284 15718 5296
rect 18322 5284 18328 5296
rect 15712 5256 18328 5284
rect 15712 5244 15718 5256
rect 18322 5244 18328 5256
rect 18380 5244 18386 5296
rect 20622 5244 20628 5296
rect 20680 5244 20686 5296
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 19889 5219 19947 5225
rect 14700 5188 15700 5216
rect 14700 5176 14706 5188
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 15672 5157 15700 5188
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5216 20591 5219
rect 20640 5216 20668 5244
rect 20806 5216 20812 5228
rect 20579 5188 20668 5216
rect 20767 5188 20812 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 13504 5120 15577 5148
rect 13504 5108 13510 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5117 15715 5151
rect 19904 5148 19932 5179
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 20254 5148 20260 5160
rect 19904 5120 20260 5148
rect 15657 5111 15715 5117
rect 15580 5012 15608 5111
rect 20254 5108 20260 5120
rect 20312 5148 20318 5160
rect 20622 5148 20628 5160
rect 20312 5120 20628 5148
rect 20312 5108 20318 5120
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 20346 5080 20352 5092
rect 20307 5052 20352 5080
rect 20346 5040 20352 5052
rect 20404 5040 20410 5092
rect 20993 5083 21051 5089
rect 20993 5049 21005 5083
rect 21039 5080 21051 5083
rect 22186 5080 22192 5092
rect 21039 5052 22192 5080
rect 21039 5049 21051 5052
rect 20993 5043 21051 5049
rect 22186 5040 22192 5052
rect 22244 5040 22250 5092
rect 16117 5015 16175 5021
rect 16117 5012 16129 5015
rect 15580 4984 16129 5012
rect 16117 4981 16129 4984
rect 16163 5012 16175 5015
rect 18230 5012 18236 5024
rect 16163 4984 18236 5012
rect 16163 4981 16175 4984
rect 16117 4975 16175 4981
rect 18230 4972 18236 4984
rect 18288 5012 18294 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18288 4984 18613 5012
rect 18288 4972 18294 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 20070 5012 20076 5024
rect 20031 4984 20076 5012
rect 18601 4975 18659 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 15436 4780 18276 4808
rect 15436 4768 15442 4780
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4641 18199 4675
rect 18248 4672 18276 4780
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 19889 4811 19947 4817
rect 19889 4808 19901 4811
rect 19760 4780 19901 4808
rect 19760 4768 19766 4780
rect 19889 4777 19901 4780
rect 19935 4777 19947 4811
rect 19889 4771 19947 4777
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20496 4780 20637 4808
rect 20496 4768 20502 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 18322 4700 18328 4752
rect 18380 4740 18386 4752
rect 20165 4743 20223 4749
rect 20165 4740 20177 4743
rect 18380 4712 20177 4740
rect 18380 4700 18386 4712
rect 20165 4709 20177 4712
rect 20211 4709 20223 4743
rect 20165 4703 20223 4709
rect 18248 4644 19840 4672
rect 18141 4635 18199 4641
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 18156 4604 18184 4635
rect 19242 4604 19248 4616
rect 16448 4576 18184 4604
rect 19203 4576 19248 4604
rect 16448 4564 16454 4576
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19444 4576 19717 4604
rect 17957 4539 18015 4545
rect 17957 4505 17969 4539
rect 18003 4536 18015 4539
rect 18601 4539 18659 4545
rect 18601 4536 18613 4539
rect 18003 4508 18613 4536
rect 18003 4505 18015 4508
rect 17957 4499 18015 4505
rect 18601 4505 18613 4508
rect 18647 4505 18659 4539
rect 18601 4499 18659 4505
rect 17034 4428 17040 4480
rect 17092 4468 17098 4480
rect 17589 4471 17647 4477
rect 17589 4468 17601 4471
rect 17092 4440 17601 4468
rect 17092 4428 17098 4440
rect 17589 4437 17601 4440
rect 17635 4437 17647 4471
rect 17589 4431 17647 4437
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18322 4468 18328 4480
rect 18095 4440 18328 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 19444 4477 19472 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19812 4536 19840 4644
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 20128 4644 20852 4672
rect 20128 4632 20134 4644
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20824 4613 20852 4644
rect 20809 4607 20867 4613
rect 20809 4573 20821 4607
rect 20855 4573 20867 4607
rect 20809 4567 20867 4573
rect 21085 4539 21143 4545
rect 21085 4536 21097 4539
rect 19812 4508 21097 4536
rect 21085 4505 21097 4508
rect 21131 4505 21143 4539
rect 21085 4499 21143 4505
rect 21269 4539 21327 4545
rect 21269 4505 21281 4539
rect 21315 4536 21327 4539
rect 21358 4536 21364 4548
rect 21315 4508 21364 4536
rect 21315 4505 21327 4508
rect 21269 4499 21327 4505
rect 21358 4496 21364 4508
rect 21416 4496 21422 4548
rect 19429 4471 19487 4477
rect 19429 4437 19441 4471
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 15194 4264 15200 4276
rect 15155 4236 15200 4264
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 17034 4264 17040 4276
rect 16995 4236 17040 4264
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 20254 4264 20260 4276
rect 20215 4236 20260 4264
rect 20254 4224 20260 4236
rect 20312 4224 20318 4276
rect 20530 4224 20536 4276
rect 20588 4264 20594 4276
rect 20625 4267 20683 4273
rect 20625 4264 20637 4267
rect 20588 4236 20637 4264
rect 20588 4224 20594 4236
rect 20625 4233 20637 4236
rect 20671 4233 20683 4267
rect 21358 4264 21364 4276
rect 20625 4227 20683 4233
rect 21100 4236 21364 4264
rect 21100 4196 21128 4236
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 21266 4196 21272 4208
rect 19904 4168 21128 4196
rect 21227 4168 21272 4196
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 14476 4100 15117 4128
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 14476 4069 14504 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 16390 4128 16396 4140
rect 15105 4091 15163 4097
rect 15764 4100 16396 4128
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 6788 4032 14473 4060
rect 6788 4020 6794 4032
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4060 15071 4063
rect 15764 4060 15792 4100
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 19904 4137 19932 4168
rect 21266 4156 21272 4168
rect 21324 4156 21330 4208
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 15059 4032 15792 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 15838 4020 15844 4072
rect 15896 4060 15902 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 15896 4032 16773 4060
rect 15896 4020 15902 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 16945 4063 17003 4069
rect 16945 4029 16957 4063
rect 16991 4029 17003 4063
rect 16945 4023 17003 4029
rect 15565 3995 15623 4001
rect 15565 3961 15577 3995
rect 15611 3992 15623 3995
rect 16960 3992 16988 4023
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 21085 4063 21143 4069
rect 21085 4060 21097 4063
rect 18288 4032 21097 4060
rect 18288 4020 18294 4032
rect 21085 4029 21097 4032
rect 21131 4029 21143 4063
rect 21085 4023 21143 4029
rect 15611 3964 16988 3992
rect 17405 3995 17463 4001
rect 15611 3961 15623 3964
rect 15565 3955 15623 3961
rect 17405 3961 17417 3995
rect 17451 3992 17463 3995
rect 19242 3992 19248 4004
rect 17451 3964 19248 3992
rect 17451 3961 17463 3964
rect 17405 3955 17463 3961
rect 19242 3952 19248 3964
rect 19300 3952 19306 4004
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 20162 3720 20168 3732
rect 20123 3692 20168 3720
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 20441 3723 20499 3729
rect 20441 3720 20453 3723
rect 20404 3692 20453 3720
rect 20404 3680 20410 3692
rect 20441 3689 20453 3692
rect 20487 3689 20499 3723
rect 20441 3683 20499 3689
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 21085 3655 21143 3661
rect 21085 3652 21097 3655
rect 15344 3624 21097 3652
rect 15344 3612 15350 3624
rect 21085 3621 21097 3624
rect 21131 3621 21143 3655
rect 21085 3615 21143 3621
rect 19797 3451 19855 3457
rect 19797 3417 19809 3451
rect 19843 3448 19855 3451
rect 21266 3448 21272 3460
rect 19843 3420 21272 3448
rect 19843 3417 19855 3420
rect 19797 3411 19855 3417
rect 21266 3408 21272 3420
rect 21324 3408 21330 3460
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 21177 3179 21235 3185
rect 21177 3176 21189 3179
rect 19576 3148 21189 3176
rect 19576 3136 19582 3148
rect 21177 3145 21189 3148
rect 21223 3145 21235 3179
rect 21177 3139 21235 3145
rect 19337 3111 19395 3117
rect 19337 3077 19349 3111
rect 19383 3108 19395 3111
rect 20622 3108 20628 3120
rect 19383 3080 20628 3108
rect 19383 3077 19395 3080
rect 19337 3071 19395 3077
rect 20622 3068 20628 3080
rect 20680 3108 20686 3120
rect 20717 3111 20775 3117
rect 20717 3108 20729 3111
rect 20680 3080 20729 3108
rect 20680 3068 20686 3080
rect 20717 3077 20729 3080
rect 20763 3077 20775 3111
rect 20717 3071 20775 3077
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 20165 3043 20223 3049
rect 20165 3040 20177 3043
rect 19751 3012 20177 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 20165 3009 20177 3012
rect 20211 3040 20223 3043
rect 20254 3040 20260 3052
rect 20211 3012 20260 3040
rect 20211 3009 20223 3012
rect 20165 3003 20223 3009
rect 20254 3000 20260 3012
rect 20312 3000 20318 3052
rect 21266 3040 21272 3052
rect 21227 3012 21272 3040
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 18969 2975 19027 2981
rect 18969 2941 18981 2975
rect 19015 2972 19027 2975
rect 21284 2972 21312 3000
rect 19015 2944 21312 2972
rect 19015 2941 19027 2944
rect 18969 2935 19027 2941
rect 17954 2864 17960 2916
rect 18012 2904 18018 2916
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 18012 2876 19993 2904
rect 18012 2864 18018 2876
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 20625 2839 20683 2845
rect 20625 2836 20637 2839
rect 15068 2808 20637 2836
rect 15068 2796 15074 2808
rect 20625 2805 20637 2808
rect 20671 2805 20683 2839
rect 20625 2799 20683 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 18874 2524 18880 2576
rect 18932 2564 18938 2576
rect 19981 2567 20039 2573
rect 19981 2564 19993 2567
rect 18932 2536 19993 2564
rect 18932 2524 18938 2536
rect 19981 2533 19993 2536
rect 20027 2533 20039 2567
rect 19981 2527 20039 2533
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 15252 2468 20821 2496
rect 15252 2456 15258 2468
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 20809 2459 20867 2465
rect 19337 2431 19395 2437
rect 19337 2397 19349 2431
rect 19383 2428 19395 2431
rect 20530 2428 20536 2440
rect 19383 2400 20536 2428
rect 19383 2397 19395 2400
rect 19337 2391 19395 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 19705 2363 19763 2369
rect 19705 2329 19717 2363
rect 19751 2360 19763 2363
rect 20162 2360 20168 2372
rect 19751 2332 20168 2360
rect 19751 2329 19763 2332
rect 19705 2323 19763 2329
rect 20162 2320 20168 2332
rect 20220 2320 20226 2372
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 5632 20544 5684 20596
rect 388 20476 440 20528
rect 1400 20476 1452 20528
rect 2044 20408 2096 20460
rect 2596 20408 2648 20460
rect 3148 20408 3200 20460
rect 4252 20408 4304 20460
rect 4804 20408 4856 20460
rect 5264 20408 5316 20460
rect 5540 20476 5592 20528
rect 5908 20476 5960 20528
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 6460 20408 6512 20460
rect 6644 20408 6696 20460
rect 6828 20408 6880 20460
rect 10416 20544 10468 20596
rect 11980 20587 12032 20596
rect 11980 20553 11989 20587
rect 11989 20553 12023 20587
rect 12023 20553 12032 20587
rect 11980 20544 12032 20553
rect 12532 20544 12584 20596
rect 13084 20544 13136 20596
rect 14740 20544 14792 20596
rect 15384 20544 15436 20596
rect 15936 20544 15988 20596
rect 17500 20544 17552 20596
rect 19340 20544 19392 20596
rect 20260 20544 20312 20596
rect 7564 20476 7616 20528
rect 9220 20476 9272 20528
rect 7104 20408 7156 20460
rect 8024 20408 8076 20460
rect 8208 20408 8260 20460
rect 9496 20408 9548 20460
rect 9772 20408 9824 20460
rect 10324 20408 10376 20460
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 10876 20408 10928 20460
rect 11060 20408 11112 20460
rect 11244 20408 11296 20460
rect 6828 20272 6880 20324
rect 7472 20272 7524 20324
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 4620 20247 4672 20256
rect 4620 20213 4629 20247
rect 4629 20213 4663 20247
rect 4663 20213 4672 20247
rect 4620 20204 4672 20213
rect 5724 20204 5776 20256
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 6736 20247 6788 20256
rect 5816 20204 5868 20213
rect 6736 20213 6745 20247
rect 6745 20213 6779 20247
rect 6779 20213 6788 20247
rect 6736 20204 6788 20213
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 7656 20247 7708 20256
rect 7656 20213 7665 20247
rect 7665 20213 7699 20247
rect 7699 20213 7708 20247
rect 7656 20204 7708 20213
rect 7748 20204 7800 20256
rect 9404 20340 9456 20392
rect 12532 20408 12584 20460
rect 12716 20408 12768 20460
rect 14648 20451 14700 20460
rect 12992 20383 13044 20392
rect 9128 20272 9180 20324
rect 12992 20349 13001 20383
rect 13001 20349 13035 20383
rect 13035 20349 13044 20383
rect 12992 20340 13044 20349
rect 13544 20340 13596 20392
rect 9680 20315 9732 20324
rect 9680 20281 9689 20315
rect 9689 20281 9723 20315
rect 9723 20281 9732 20315
rect 9680 20272 9732 20281
rect 13084 20272 13136 20324
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 16212 20408 16264 20460
rect 17040 20408 17092 20460
rect 17592 20408 17644 20460
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 19616 20476 19668 20528
rect 19892 20408 19944 20460
rect 21180 20476 21232 20528
rect 20904 20451 20956 20460
rect 15292 20340 15344 20392
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 20996 20340 21048 20392
rect 9312 20204 9364 20256
rect 10508 20247 10560 20256
rect 10508 20213 10517 20247
rect 10517 20213 10551 20247
rect 10551 20213 10560 20247
rect 10508 20204 10560 20213
rect 12164 20204 12216 20256
rect 12440 20204 12492 20256
rect 14188 20272 14240 20324
rect 16948 20272 17000 20324
rect 18144 20272 18196 20324
rect 19524 20272 19576 20324
rect 19708 20272 19760 20324
rect 13452 20204 13504 20256
rect 16580 20204 16632 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 2596 20043 2648 20052
rect 2596 20009 2605 20043
rect 2605 20009 2639 20043
rect 2639 20009 2648 20043
rect 2596 20000 2648 20009
rect 3148 20000 3200 20052
rect 3424 20043 3476 20052
rect 3424 20009 3433 20043
rect 3433 20009 3467 20043
rect 3467 20009 3476 20043
rect 3424 20000 3476 20009
rect 4804 20000 4856 20052
rect 6000 20000 6052 20052
rect 9128 20043 9180 20052
rect 5540 19932 5592 19984
rect 8852 19932 8904 19984
rect 6828 19907 6880 19916
rect 1492 19796 1544 19848
rect 3424 19796 3476 19848
rect 6828 19873 6837 19907
rect 6837 19873 6871 19907
rect 6871 19873 6880 19907
rect 6828 19864 6880 19873
rect 8024 19864 8076 19916
rect 9128 20009 9137 20043
rect 9137 20009 9171 20043
rect 9171 20009 9180 20043
rect 9128 20000 9180 20009
rect 9404 20043 9456 20052
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 13544 20043 13596 20052
rect 9036 19932 9088 19984
rect 9864 19975 9916 19984
rect 9864 19941 9873 19975
rect 9873 19941 9907 19975
rect 9907 19941 9916 19975
rect 9864 19932 9916 19941
rect 7012 19728 7064 19780
rect 1768 19703 1820 19712
rect 1768 19669 1777 19703
rect 1777 19669 1811 19703
rect 1811 19669 1820 19703
rect 1768 19660 1820 19669
rect 3976 19703 4028 19712
rect 3976 19669 3985 19703
rect 3985 19669 4019 19703
rect 4019 19669 4028 19703
rect 3976 19660 4028 19669
rect 5908 19703 5960 19712
rect 5908 19669 5917 19703
rect 5917 19669 5951 19703
rect 5951 19669 5960 19703
rect 5908 19660 5960 19669
rect 7380 19728 7432 19780
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 8484 19660 8536 19712
rect 8668 19796 8720 19848
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 10968 19839 11020 19848
rect 10968 19805 10986 19839
rect 10986 19805 11020 19839
rect 11244 19839 11296 19848
rect 10968 19796 11020 19805
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 13820 20000 13872 20052
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 17868 20000 17920 20052
rect 18604 20000 18656 20052
rect 15292 19975 15344 19984
rect 12716 19864 12768 19916
rect 12624 19796 12676 19848
rect 11704 19728 11756 19780
rect 12440 19728 12492 19780
rect 11152 19660 11204 19712
rect 15292 19941 15301 19975
rect 15301 19941 15335 19975
rect 15335 19941 15344 19975
rect 15292 19932 15344 19941
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 13452 19864 13504 19916
rect 14464 19796 14516 19848
rect 14832 19839 14884 19848
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 17224 19864 17276 19916
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 17132 19796 17184 19848
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 18420 19907 18472 19916
rect 18420 19873 18429 19907
rect 18429 19873 18463 19907
rect 18463 19873 18472 19907
rect 18604 19907 18656 19916
rect 18420 19864 18472 19873
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19800 19864 19852 19916
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 16396 19728 16448 19780
rect 13176 19703 13228 19712
rect 13176 19669 13185 19703
rect 13185 19669 13219 19703
rect 13219 19669 13228 19703
rect 13176 19660 13228 19669
rect 15844 19703 15896 19712
rect 15844 19669 15853 19703
rect 15853 19669 15887 19703
rect 15887 19669 15896 19703
rect 15844 19660 15896 19669
rect 17408 19660 17460 19712
rect 17776 19660 17828 19712
rect 18236 19660 18288 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 1492 19456 1544 19508
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 5908 19456 5960 19508
rect 7104 19456 7156 19508
rect 7932 19499 7984 19508
rect 7932 19465 7941 19499
rect 7941 19465 7975 19499
rect 7975 19465 7984 19499
rect 7932 19456 7984 19465
rect 8024 19456 8076 19508
rect 4712 19363 4764 19372
rect 940 19252 992 19304
rect 4712 19329 4721 19363
rect 4721 19329 4755 19363
rect 4755 19329 4764 19363
rect 4712 19320 4764 19329
rect 6644 19388 6696 19440
rect 8208 19388 8260 19440
rect 6920 19320 6972 19372
rect 8300 19320 8352 19372
rect 9588 19456 9640 19508
rect 11704 19456 11756 19508
rect 11796 19456 11848 19508
rect 17224 19456 17276 19508
rect 19616 19499 19668 19508
rect 9680 19320 9732 19372
rect 11244 19388 11296 19440
rect 11888 19388 11940 19440
rect 12624 19388 12676 19440
rect 16028 19388 16080 19440
rect 9864 19320 9916 19372
rect 11152 19320 11204 19372
rect 12716 19320 12768 19372
rect 12992 19320 13044 19372
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 8208 19252 8260 19304
rect 9772 19184 9824 19236
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 7380 19116 7432 19168
rect 12072 19184 12124 19236
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 18512 19320 18564 19372
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19064 19320 19116 19372
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 20628 19456 20680 19508
rect 18052 19252 18104 19304
rect 17960 19184 18012 19236
rect 19156 19252 19208 19304
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 20812 19320 20864 19372
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 12532 19159 12584 19168
rect 12532 19125 12541 19159
rect 12541 19125 12575 19159
rect 12575 19125 12584 19159
rect 12532 19116 12584 19125
rect 14372 19116 14424 19168
rect 17224 19116 17276 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1400 18955 1452 18964
rect 1400 18921 1409 18955
rect 1409 18921 1443 18955
rect 1443 18921 1452 18955
rect 1400 18912 1452 18921
rect 7012 18955 7064 18964
rect 7012 18921 7021 18955
rect 7021 18921 7055 18955
rect 7055 18921 7064 18955
rect 7012 18912 7064 18921
rect 9220 18912 9272 18964
rect 10692 18912 10744 18964
rect 11060 18912 11112 18964
rect 18052 18955 18104 18964
rect 18052 18921 18061 18955
rect 18061 18921 18095 18955
rect 18095 18921 18104 18955
rect 18052 18912 18104 18921
rect 21364 18912 21416 18964
rect 6552 18844 6604 18896
rect 5724 18776 5776 18828
rect 9404 18844 9456 18896
rect 18880 18844 18932 18896
rect 7472 18819 7524 18828
rect 7472 18785 7481 18819
rect 7481 18785 7515 18819
rect 7515 18785 7524 18819
rect 7472 18776 7524 18785
rect 7840 18572 7892 18624
rect 9404 18572 9456 18624
rect 10968 18640 11020 18692
rect 11244 18640 11296 18692
rect 13820 18708 13872 18760
rect 18696 18776 18748 18828
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 17408 18708 17460 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 11888 18572 11940 18624
rect 12072 18572 12124 18624
rect 13176 18572 13228 18624
rect 13544 18572 13596 18624
rect 16948 18572 17000 18624
rect 17868 18572 17920 18624
rect 20260 18640 20312 18692
rect 21548 18640 21600 18692
rect 21088 18572 21140 18624
rect 21364 18572 21416 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 7564 18368 7616 18420
rect 10508 18368 10560 18420
rect 18972 18368 19024 18420
rect 6644 18300 6696 18352
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 8208 18232 8260 18284
rect 6552 18164 6604 18216
rect 11796 18300 11848 18352
rect 12716 18300 12768 18352
rect 16856 18300 16908 18352
rect 17224 18300 17276 18352
rect 9680 18232 9732 18284
rect 5540 18096 5592 18148
rect 8392 18096 8444 18148
rect 8576 18028 8628 18080
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 10784 18028 10836 18080
rect 11888 18232 11940 18284
rect 15936 18207 15988 18216
rect 15936 18173 15945 18207
rect 15945 18173 15979 18207
rect 15979 18173 15988 18207
rect 15936 18164 15988 18173
rect 16948 18232 17000 18284
rect 18972 18232 19024 18284
rect 19524 18232 19576 18284
rect 19708 18232 19760 18284
rect 20444 18232 20496 18284
rect 21088 18275 21140 18284
rect 21088 18241 21097 18275
rect 21097 18241 21131 18275
rect 21131 18241 21140 18275
rect 21088 18232 21140 18241
rect 11888 18028 11940 18080
rect 14280 18028 14332 18080
rect 14372 18028 14424 18080
rect 19800 18096 19852 18148
rect 20168 18139 20220 18148
rect 20168 18105 20177 18139
rect 20177 18105 20211 18139
rect 20211 18105 20220 18139
rect 20168 18096 20220 18105
rect 17868 18028 17920 18080
rect 22468 18096 22520 18148
rect 20628 18028 20680 18080
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 4712 17824 4764 17876
rect 9772 17824 9824 17876
rect 16120 17824 16172 17876
rect 16396 17824 16448 17876
rect 17500 17867 17552 17876
rect 17500 17833 17509 17867
rect 17509 17833 17543 17867
rect 17543 17833 17552 17867
rect 17500 17824 17552 17833
rect 17960 17824 18012 17876
rect 6644 17731 6696 17740
rect 6644 17697 6653 17731
rect 6653 17697 6687 17731
rect 6687 17697 6696 17731
rect 6644 17688 6696 17697
rect 16856 17756 16908 17808
rect 7748 17688 7800 17740
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 5540 17552 5592 17604
rect 9128 17688 9180 17740
rect 17868 17688 17920 17740
rect 19340 17688 19392 17740
rect 15936 17620 15988 17672
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 8576 17484 8628 17536
rect 19800 17620 19852 17672
rect 18604 17595 18656 17604
rect 18604 17561 18622 17595
rect 18622 17561 18656 17595
rect 18604 17552 18656 17561
rect 17500 17484 17552 17536
rect 19616 17484 19668 17536
rect 20628 17552 20680 17604
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 5540 17323 5592 17332
rect 5540 17289 5549 17323
rect 5549 17289 5583 17323
rect 5583 17289 5592 17323
rect 5540 17280 5592 17289
rect 8392 17280 8444 17332
rect 16028 17323 16080 17332
rect 16028 17289 16037 17323
rect 16037 17289 16071 17323
rect 16071 17289 16080 17323
rect 16028 17280 16080 17289
rect 16948 17280 17000 17332
rect 19340 17280 19392 17332
rect 21088 17280 21140 17332
rect 4804 17212 4856 17264
rect 10876 17187 10928 17196
rect 10876 17153 10894 17187
rect 10894 17153 10928 17187
rect 10876 17144 10928 17153
rect 4160 17008 4212 17060
rect 8024 17008 8076 17060
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11888 16940 11940 16992
rect 14280 17212 14332 17264
rect 13820 17144 13872 17196
rect 15844 17144 15896 17196
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 17684 17008 17736 17060
rect 19616 17144 19668 17196
rect 20076 17144 20128 17196
rect 20720 17144 20772 17196
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 19524 16940 19576 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20536 16940 20588 16992
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 4620 16736 4672 16788
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 5816 16668 5868 16720
rect 5540 16532 5592 16584
rect 18604 16736 18656 16788
rect 20628 16736 20680 16788
rect 9772 16668 9824 16720
rect 18788 16711 18840 16720
rect 18788 16677 18797 16711
rect 18797 16677 18831 16711
rect 18831 16677 18840 16711
rect 18788 16668 18840 16677
rect 7932 16643 7984 16652
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 7840 16464 7892 16516
rect 9772 16532 9824 16584
rect 14372 16600 14424 16652
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 18144 16575 18196 16584
rect 18144 16541 18153 16575
rect 18153 16541 18187 16575
rect 18187 16541 18196 16575
rect 18144 16532 18196 16541
rect 11704 16464 11756 16516
rect 12256 16464 12308 16516
rect 21364 16532 21416 16584
rect 5264 16396 5316 16448
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 6000 16396 6052 16405
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 7288 16396 7340 16448
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 8392 16396 8444 16448
rect 11244 16396 11296 16448
rect 13820 16396 13872 16448
rect 19524 16396 19576 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 7288 16235 7340 16244
rect 7288 16201 7297 16235
rect 7297 16201 7331 16235
rect 7331 16201 7340 16235
rect 7288 16192 7340 16201
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 12256 16192 12308 16244
rect 12992 16124 13044 16176
rect 14372 16192 14424 16244
rect 15292 16124 15344 16176
rect 20076 16192 20128 16244
rect 20628 16192 20680 16244
rect 20720 16124 20772 16176
rect 5448 16056 5500 16108
rect 10876 15988 10928 16040
rect 11888 15988 11940 16040
rect 17960 16056 18012 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 19800 16056 19852 16108
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20352 15988 20404 16040
rect 6000 15852 6052 15904
rect 9128 15852 9180 15904
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 11888 15852 11940 15904
rect 15292 15852 15344 15904
rect 17684 15895 17736 15904
rect 17684 15861 17693 15895
rect 17693 15861 17727 15895
rect 17727 15861 17736 15895
rect 17684 15852 17736 15861
rect 18236 15852 18288 15904
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 7012 15648 7064 15700
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 7656 15512 7708 15564
rect 12256 15648 12308 15700
rect 19064 15648 19116 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20444 15648 20496 15700
rect 17684 15512 17736 15564
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 11520 15444 11572 15496
rect 12348 15444 12400 15496
rect 18236 15487 18288 15496
rect 10048 15419 10100 15428
rect 10048 15385 10082 15419
rect 10082 15385 10100 15419
rect 10048 15376 10100 15385
rect 12808 15376 12860 15428
rect 16396 15376 16448 15428
rect 8392 15308 8444 15360
rect 11060 15308 11112 15360
rect 15844 15308 15896 15360
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 22192 15444 22244 15496
rect 20720 15376 20772 15428
rect 17868 15308 17920 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 5632 15104 5684 15156
rect 17132 15147 17184 15156
rect 7932 15036 7984 15088
rect 9588 15036 9640 15088
rect 12348 15036 12400 15088
rect 9772 14968 9824 15020
rect 12256 14968 12308 15020
rect 7104 14900 7156 14952
rect 10876 14832 10928 14884
rect 11704 14832 11756 14884
rect 11244 14764 11296 14816
rect 14280 14764 14332 14816
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 20168 15104 20220 15156
rect 20536 15147 20588 15156
rect 20536 15113 20545 15147
rect 20545 15113 20579 15147
rect 20579 15113 20588 15147
rect 20536 15104 20588 15113
rect 17500 14968 17552 15020
rect 22100 14968 22152 15020
rect 20812 14832 20864 14884
rect 19800 14764 19852 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 16672 14560 16724 14612
rect 17500 14560 17552 14612
rect 19524 14560 19576 14612
rect 20628 14560 20680 14612
rect 11060 14424 11112 14476
rect 7564 14356 7616 14408
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 15844 14288 15896 14340
rect 17868 14356 17920 14408
rect 20076 14356 20128 14408
rect 21640 14356 21692 14408
rect 17040 14288 17092 14340
rect 18788 14220 18840 14272
rect 19616 14220 19668 14272
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 7564 14016 7616 14068
rect 8300 14059 8352 14068
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9588 14016 9640 14025
rect 11244 14016 11296 14068
rect 11612 14016 11664 14068
rect 12808 14059 12860 14068
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 11060 13948 11112 14000
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 11796 13948 11848 14000
rect 14648 13948 14700 14000
rect 19892 13948 19944 14000
rect 19524 13923 19576 13932
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 20812 14016 20864 14068
rect 21180 14059 21232 14068
rect 21180 14025 21189 14059
rect 21189 14025 21223 14059
rect 21223 14025 21232 14059
rect 21180 14016 21232 14025
rect 20628 13880 20680 13932
rect 21456 13880 21508 13932
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 14280 13812 14332 13864
rect 12808 13744 12860 13796
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 15016 13676 15068 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 7380 13472 7432 13524
rect 3976 13336 4028 13388
rect 10048 13472 10100 13524
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 16396 13515 16448 13524
rect 8392 13200 8444 13252
rect 9772 13200 9824 13252
rect 11888 13200 11940 13252
rect 11980 13132 12032 13184
rect 12072 13132 12124 13184
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 17868 13472 17920 13524
rect 17040 13404 17092 13456
rect 19524 13472 19576 13524
rect 20260 13472 20312 13524
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 15292 13311 15344 13320
rect 15292 13277 15326 13311
rect 15326 13277 15344 13311
rect 15292 13268 15344 13277
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 20996 13268 21048 13320
rect 21180 13268 21232 13320
rect 14832 13200 14884 13252
rect 16488 13132 16540 13184
rect 17040 13200 17092 13252
rect 18052 13200 18104 13252
rect 18696 13132 18748 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 7012 12928 7064 12980
rect 7288 12928 7340 12980
rect 8024 12792 8076 12844
rect 10140 12792 10192 12844
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 11704 12928 11756 12980
rect 11980 12928 12032 12980
rect 13820 12928 13872 12980
rect 16396 12928 16448 12980
rect 15016 12860 15068 12912
rect 19524 12928 19576 12980
rect 19984 12928 20036 12980
rect 21088 12928 21140 12980
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 14280 12835 14332 12844
rect 14280 12801 14314 12835
rect 14314 12801 14332 12835
rect 14280 12792 14332 12801
rect 18788 12792 18840 12844
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 5540 12588 5592 12640
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 11796 12588 11848 12640
rect 13820 12588 13872 12640
rect 14924 12588 14976 12640
rect 17040 12588 17092 12640
rect 18880 12588 18932 12640
rect 21364 12588 21416 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 5540 12248 5592 12300
rect 5908 12248 5960 12300
rect 12072 12384 12124 12436
rect 20260 12427 20312 12436
rect 20260 12393 20269 12427
rect 20269 12393 20303 12427
rect 20303 12393 20312 12427
rect 20260 12384 20312 12393
rect 20904 12427 20956 12436
rect 20904 12393 20913 12427
rect 20913 12393 20947 12427
rect 20947 12393 20956 12427
rect 20904 12384 20956 12393
rect 20996 12384 21048 12436
rect 20536 12316 20588 12368
rect 10140 12248 10192 12300
rect 8208 12180 8260 12232
rect 8300 12180 8352 12232
rect 14556 12248 14608 12300
rect 5080 12087 5132 12096
rect 5080 12053 5089 12087
rect 5089 12053 5123 12087
rect 5123 12053 5132 12087
rect 5448 12087 5500 12096
rect 5080 12044 5132 12053
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 10508 12112 10560 12164
rect 8024 12044 8076 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 13912 12180 13964 12232
rect 15016 12180 15068 12232
rect 16120 12112 16172 12164
rect 11704 12044 11756 12096
rect 14280 12044 14332 12096
rect 19064 12044 19116 12096
rect 21180 12180 21232 12232
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 21548 12112 21600 12164
rect 21640 12044 21692 12096
rect 22284 12044 22336 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 5080 11840 5132 11892
rect 8668 11840 8720 11892
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 18696 11840 18748 11892
rect 18972 11840 19024 11892
rect 21548 11840 21600 11892
rect 20812 11772 20864 11824
rect 21272 11772 21324 11824
rect 21640 11772 21692 11824
rect 8208 11704 8260 11756
rect 21364 11704 21416 11756
rect 21272 11636 21324 11688
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 19524 11500 19576 11552
rect 19616 11543 19668 11552
rect 19616 11509 19625 11543
rect 19625 11509 19659 11543
rect 19659 11509 19668 11543
rect 19616 11500 19668 11509
rect 19892 11500 19944 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 13820 11296 13872 11348
rect 14556 11296 14608 11348
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 12348 11135 12400 11144
rect 11704 11092 11756 11101
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12440 11092 12492 11144
rect 20812 11228 20864 11280
rect 18788 11092 18840 11144
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 12992 11024 13044 11076
rect 15108 11024 15160 11076
rect 13728 10999 13780 11008
rect 13728 10965 13737 10999
rect 13737 10965 13771 10999
rect 13771 10965 13780 10999
rect 13728 10956 13780 10965
rect 15016 10956 15068 11008
rect 18328 11024 18380 11076
rect 19064 11024 19116 11076
rect 19800 11024 19852 11076
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 1584 10752 1636 10804
rect 8024 10616 8076 10668
rect 9772 10616 9824 10668
rect 10876 10616 10928 10668
rect 12348 10684 12400 10736
rect 8208 10548 8260 10600
rect 15108 10684 15160 10736
rect 18236 10752 18288 10804
rect 20904 10752 20956 10804
rect 13728 10616 13780 10668
rect 8300 10480 8352 10532
rect 8024 10412 8076 10464
rect 10968 10412 11020 10464
rect 12900 10548 12952 10600
rect 15108 10548 15160 10600
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 17868 10480 17920 10532
rect 19800 10616 19852 10668
rect 21272 10684 21324 10736
rect 21548 10548 21600 10600
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 14372 10412 14424 10464
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 12348 10208 12400 10260
rect 11888 10140 11940 10192
rect 15108 10208 15160 10260
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 14464 10004 14516 10056
rect 19524 10072 19576 10124
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 9956 9979 10008 9988
rect 9956 9945 9990 9979
rect 9990 9945 10008 9979
rect 9956 9936 10008 9945
rect 13820 9936 13872 9988
rect 16672 9936 16724 9988
rect 19800 9936 19852 9988
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 8300 9664 8352 9716
rect 20352 9664 20404 9716
rect 10416 9596 10468 9648
rect 18144 9596 18196 9648
rect 18420 9596 18472 9648
rect 8576 9528 8628 9580
rect 9404 9528 9456 9580
rect 13544 9528 13596 9580
rect 19800 9528 19852 9580
rect 20260 9571 20312 9580
rect 10876 9460 10928 9512
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 20996 9460 21048 9512
rect 7840 9392 7892 9444
rect 14648 9392 14700 9444
rect 19984 9392 20036 9444
rect 20444 9435 20496 9444
rect 20444 9401 20453 9435
rect 20453 9401 20487 9435
rect 20487 9401 20496 9435
rect 20444 9392 20496 9401
rect 20720 9435 20772 9444
rect 20720 9401 20729 9435
rect 20729 9401 20763 9435
rect 20763 9401 20772 9435
rect 20720 9392 20772 9401
rect 21456 9392 21508 9444
rect 10692 9324 10744 9376
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 16212 9324 16264 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 10508 9120 10560 9172
rect 8208 8984 8260 9036
rect 10968 9052 11020 9104
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 8116 8916 8168 8968
rect 20260 9120 20312 9172
rect 21088 9163 21140 9172
rect 21088 9129 21097 9163
rect 21097 9129 21131 9163
rect 21131 9129 21140 9163
rect 21088 9120 21140 9129
rect 11888 9052 11940 9104
rect 13820 8984 13872 9036
rect 7840 8780 7892 8832
rect 10416 8848 10468 8900
rect 12072 8848 12124 8900
rect 15384 8984 15436 9036
rect 19064 8984 19116 9036
rect 19800 9027 19852 9036
rect 19800 8993 19809 9027
rect 19809 8993 19843 9027
rect 19843 8993 19852 9027
rect 19800 8984 19852 8993
rect 20628 9027 20680 9036
rect 20628 8993 20637 9027
rect 20637 8993 20671 9027
rect 20671 8993 20680 9027
rect 20628 8984 20680 8993
rect 16120 8916 16172 8968
rect 17132 8916 17184 8968
rect 19248 8959 19300 8968
rect 9404 8780 9456 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 11152 8823 11204 8832
rect 10784 8780 10836 8789
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 11796 8823 11848 8832
rect 11796 8789 11805 8823
rect 11805 8789 11839 8823
rect 11839 8789 11848 8823
rect 11796 8780 11848 8789
rect 12256 8780 12308 8832
rect 13176 8780 13228 8832
rect 13544 8780 13596 8832
rect 14464 8780 14516 8832
rect 14924 8780 14976 8832
rect 16304 8848 16356 8900
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 20536 8916 20588 8968
rect 22100 8848 22152 8900
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 19064 8780 19116 8832
rect 20076 8823 20128 8832
rect 20076 8789 20085 8823
rect 20085 8789 20119 8823
rect 20119 8789 20128 8823
rect 20076 8780 20128 8789
rect 20536 8823 20588 8832
rect 20536 8789 20545 8823
rect 20545 8789 20579 8823
rect 20579 8789 20588 8823
rect 20536 8780 20588 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 10784 8576 10836 8628
rect 11152 8576 11204 8628
rect 12256 8619 12308 8628
rect 2320 8372 2372 8424
rect 11704 8508 11756 8560
rect 12256 8585 12265 8619
rect 12265 8585 12299 8619
rect 12299 8585 12308 8619
rect 12256 8576 12308 8585
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 14648 8576 14700 8628
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 16304 8576 16356 8628
rect 17132 8619 17184 8628
rect 11244 8440 11296 8492
rect 14464 8508 14516 8560
rect 15292 8508 15344 8560
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 18144 8576 18196 8628
rect 19892 8576 19944 8628
rect 20536 8576 20588 8628
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 10692 8372 10744 8424
rect 10876 8415 10928 8424
rect 10876 8381 10885 8415
rect 10885 8381 10919 8415
rect 10919 8381 10928 8415
rect 10876 8372 10928 8381
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 8024 8304 8076 8356
rect 12440 8372 12492 8424
rect 16212 8440 16264 8492
rect 15200 8304 15252 8356
rect 15476 8372 15528 8424
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 19800 8440 19852 8492
rect 20352 8483 20404 8492
rect 20352 8449 20361 8483
rect 20361 8449 20395 8483
rect 20395 8449 20404 8483
rect 20352 8440 20404 8449
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 17408 8372 17460 8424
rect 18328 8372 18380 8424
rect 17960 8304 18012 8356
rect 18880 8304 18932 8356
rect 20904 8304 20956 8356
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 20720 8236 20772 8288
rect 21640 8236 21692 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 17500 8032 17552 8084
rect 20352 8032 20404 8084
rect 20996 8032 21048 8084
rect 11060 7964 11112 8016
rect 12072 8007 12124 8016
rect 12072 7973 12081 8007
rect 12081 7973 12115 8007
rect 12115 7973 12124 8007
rect 12072 7964 12124 7973
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 20536 7964 20588 8016
rect 20720 8007 20772 8016
rect 20720 7973 20729 8007
rect 20729 7973 20763 8007
rect 20763 7973 20772 8007
rect 20720 7964 20772 7973
rect 21180 7964 21232 8016
rect 22284 7964 22336 8016
rect 13820 7828 13872 7880
rect 15200 7828 15252 7880
rect 17868 7896 17920 7948
rect 19248 7896 19300 7948
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 15016 7692 15068 7744
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 20904 7871 20956 7880
rect 19892 7803 19944 7812
rect 19892 7769 19901 7803
rect 19901 7769 19935 7803
rect 19935 7769 19944 7803
rect 19892 7760 19944 7769
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 20996 7828 21048 7880
rect 21180 7828 21232 7880
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 20996 7692 21048 7744
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 21364 7692 21416 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 20076 7488 20128 7540
rect 21088 7488 21140 7540
rect 11888 7420 11940 7472
rect 2872 7352 2924 7404
rect 21456 7352 21508 7404
rect 21548 7284 21600 7336
rect 14280 7216 14332 7268
rect 14924 7216 14976 7268
rect 20168 7216 20220 7268
rect 13636 7148 13688 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15936 7148 15988 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 13636 6808 13688 6860
rect 13728 6740 13780 6792
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 14924 6808 14976 6860
rect 17040 6808 17092 6860
rect 17776 6808 17828 6860
rect 19616 6808 19668 6860
rect 19984 6808 20036 6860
rect 21364 6851 21416 6860
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 9128 6672 9180 6724
rect 13820 6604 13872 6656
rect 13912 6604 13964 6656
rect 14832 6672 14884 6724
rect 15200 6604 15252 6656
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 17500 6672 17552 6724
rect 15752 6604 15804 6613
rect 17224 6604 17276 6656
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 17684 6604 17736 6656
rect 18052 6604 18104 6656
rect 20260 6604 20312 6656
rect 20628 6604 20680 6656
rect 20720 6604 20772 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 14832 6400 14884 6452
rect 15752 6443 15804 6452
rect 15752 6409 15761 6443
rect 15761 6409 15795 6443
rect 15795 6409 15804 6443
rect 15752 6400 15804 6409
rect 15936 6400 15988 6452
rect 1768 6332 1820 6384
rect 13912 6332 13964 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 15200 6332 15252 6384
rect 11888 6264 11940 6273
rect 15108 6264 15160 6316
rect 17500 6400 17552 6452
rect 17684 6443 17736 6452
rect 17684 6409 17693 6443
rect 17693 6409 17727 6443
rect 17727 6409 17736 6443
rect 17684 6400 17736 6409
rect 19524 6443 19576 6452
rect 19524 6409 19533 6443
rect 19533 6409 19567 6443
rect 19567 6409 19576 6443
rect 19524 6400 19576 6409
rect 20260 6443 20312 6452
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 20628 6443 20680 6452
rect 20628 6409 20637 6443
rect 20637 6409 20671 6443
rect 20671 6409 20680 6443
rect 20628 6400 20680 6409
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 17316 6332 17368 6384
rect 12900 6239 12952 6248
rect 9956 6128 10008 6180
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 14372 6239 14424 6248
rect 12992 6128 13044 6180
rect 13728 6171 13780 6180
rect 13728 6137 13737 6171
rect 13737 6137 13771 6171
rect 13771 6137 13780 6171
rect 13728 6128 13780 6137
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 14648 6128 14700 6180
rect 12348 6060 12400 6112
rect 18880 6307 18932 6316
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 18880 6273 18889 6307
rect 18889 6273 18923 6307
rect 18923 6273 18932 6307
rect 18880 6264 18932 6273
rect 19892 6332 19944 6384
rect 20536 6332 20588 6384
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 19524 6128 19576 6180
rect 14924 6060 14976 6112
rect 18144 6060 18196 6112
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 20812 6060 20864 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 17868 5856 17920 5908
rect 18144 5856 18196 5908
rect 18788 5899 18840 5908
rect 18788 5865 18797 5899
rect 18797 5865 18831 5899
rect 18831 5865 18840 5899
rect 18788 5856 18840 5865
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 20536 5856 20588 5908
rect 17592 5788 17644 5840
rect 20720 5831 20772 5840
rect 20720 5797 20729 5831
rect 20729 5797 20763 5831
rect 20763 5797 20772 5831
rect 20720 5788 20772 5797
rect 12900 5720 12952 5772
rect 18236 5720 18288 5772
rect 19064 5720 19116 5772
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 15568 5559 15620 5568
rect 15568 5525 15577 5559
rect 15577 5525 15611 5559
rect 15611 5525 15620 5559
rect 15568 5516 15620 5525
rect 18328 5584 18380 5636
rect 21180 5584 21232 5636
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 19524 5516 19576 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 15568 5312 15620 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 19984 5312 20036 5364
rect 20352 5312 20404 5364
rect 15660 5244 15712 5296
rect 18328 5244 18380 5296
rect 20628 5244 20680 5296
rect 14648 5176 14700 5228
rect 13452 5108 13504 5160
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 20260 5108 20312 5160
rect 20628 5108 20680 5160
rect 20352 5083 20404 5092
rect 20352 5049 20361 5083
rect 20361 5049 20395 5083
rect 20395 5049 20404 5083
rect 20352 5040 20404 5049
rect 22192 5040 22244 5092
rect 18236 4972 18288 5024
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 15384 4768 15436 4820
rect 19708 4768 19760 4820
rect 20444 4768 20496 4820
rect 18328 4700 18380 4752
rect 16396 4564 16448 4616
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 17040 4428 17092 4480
rect 18328 4428 18380 4480
rect 20076 4632 20128 4684
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 21364 4496 21416 4548
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 15200 4267 15252 4276
rect 15200 4233 15209 4267
rect 15209 4233 15243 4267
rect 15243 4233 15252 4267
rect 15200 4224 15252 4233
rect 17040 4267 17092 4276
rect 17040 4233 17049 4267
rect 17049 4233 17083 4267
rect 17083 4233 17092 4267
rect 17040 4224 17092 4233
rect 20260 4267 20312 4276
rect 20260 4233 20269 4267
rect 20269 4233 20303 4267
rect 20303 4233 20312 4267
rect 20260 4224 20312 4233
rect 20536 4224 20588 4276
rect 21364 4224 21416 4276
rect 21272 4199 21324 4208
rect 6736 4020 6788 4072
rect 16396 4088 16448 4140
rect 21272 4165 21281 4199
rect 21281 4165 21315 4199
rect 21315 4165 21324 4199
rect 21272 4156 21324 4165
rect 15844 4020 15896 4072
rect 18236 4020 18288 4072
rect 19248 3952 19300 4004
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 20168 3723 20220 3732
rect 20168 3689 20177 3723
rect 20177 3689 20211 3723
rect 20211 3689 20220 3723
rect 20168 3680 20220 3689
rect 20352 3680 20404 3732
rect 15292 3612 15344 3664
rect 21272 3451 21324 3460
rect 21272 3417 21281 3451
rect 21281 3417 21315 3451
rect 21315 3417 21324 3451
rect 21272 3408 21324 3417
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 19524 3136 19576 3188
rect 20628 3068 20680 3120
rect 20260 3000 20312 3052
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 17960 2864 18012 2916
rect 15016 2796 15068 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 18880 2524 18932 2576
rect 15200 2456 15252 2508
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 20168 2363 20220 2372
rect 20168 2329 20177 2363
rect 20177 2329 20211 2363
rect 20211 2329 20220 2363
rect 20168 2320 20220 2329
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
<< metal2 >>
rect 386 22200 442 23000
rect 938 22200 994 23000
rect 1490 22200 1546 23000
rect 2042 22200 2098 23000
rect 2594 22200 2650 23000
rect 3146 22200 3202 23000
rect 3436 22222 3648 22250
rect 400 20534 428 22200
rect 388 20528 440 20534
rect 388 20470 440 20476
rect 952 19310 980 22200
rect 1400 20528 1452 20534
rect 1400 20470 1452 20476
rect 940 19304 992 19310
rect 940 19246 992 19252
rect 1412 18970 1440 20470
rect 1504 19854 1532 22200
rect 2056 20466 2084 22200
rect 2608 20466 2636 22200
rect 3160 20466 3188 22200
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 2056 20058 2084 20402
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 1504 19514 1532 19790
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1596 10810 1624 19110
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1780 6390 1808 19654
rect 2332 8430 2360 20198
rect 2608 20058 2636 20402
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2884 7410 2912 20198
rect 3160 20058 3188 20402
rect 3436 20058 3464 22222
rect 3620 22114 3648 22222
rect 3698 22200 3754 23000
rect 4250 22200 4306 23000
rect 4802 22200 4858 23000
rect 5354 22200 5410 23000
rect 5906 22200 5962 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8312 22222 8616 22250
rect 3712 22114 3740 22200
rect 3620 22086 3740 22114
rect 4264 20466 4292 22200
rect 4816 20466 4844 22200
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 5264 20460 5316 20466
rect 5368 20448 5396 22200
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5316 20420 5396 20448
rect 5264 20402 5316 20408
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3436 19854 3464 19994
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3988 13394 4016 19654
rect 4172 17066 4200 20198
rect 4264 19310 4292 20402
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4632 16794 4660 20198
rect 4816 20058 4844 20402
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 5276 19514 5304 20402
rect 5552 19990 5580 20470
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4724 17882 4752 19314
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 5184 17678 5212 18158
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5552 17610 5580 18090
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4816 16658 4844 17206
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 5552 16590 5580 17274
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5644 16538 5672 20538
rect 5920 20534 5948 22200
rect 6472 20890 6500 22200
rect 6472 20862 6592 20890
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 5908 20528 5960 20534
rect 5908 20470 5960 20476
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6460 20460 6512 20466
rect 6564 20448 6592 20862
rect 6512 20420 6592 20448
rect 6644 20460 6696 20466
rect 6460 20402 6512 20408
rect 6644 20402 6696 20408
rect 6828 20460 6880 20466
rect 7024 20448 7052 22200
rect 7576 20534 7604 22200
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 6880 20420 7052 20448
rect 7104 20460 7156 20466
rect 6828 20402 6880 20408
rect 7104 20402 7156 20408
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5736 18834 5764 20198
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5828 16726 5856 20198
rect 6012 20058 6040 20402
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5920 19514 5948 19654
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 6656 19446 6684 20402
rect 6828 20324 6880 20330
rect 6828 20266 6880 20272
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6564 18222 6592 18838
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6656 17746 6684 18294
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 5644 16510 5948 16538
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5276 16250 5304 16390
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15570 5488 16050
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5644 15162 5672 16390
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 5552 12306 5580 12582
rect 5920 12306 5948 16510
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 6012 15910 6040 16390
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5092 11898 5120 12038
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 5460 9081 5488 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 5446 9072 5502 9081
rect 5446 9007 5502 9016
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5817 1440 6258
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6748 4078 6776 20198
rect 6840 19922 6868 20266
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6918 19816 6974 19825
rect 6918 19751 6974 19760
rect 7012 19780 7064 19786
rect 6932 19378 6960 19751
rect 7012 19722 7064 19728
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7024 18970 7052 19722
rect 7116 19514 7144 20402
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 15706 7052 16390
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 14074 7144 14894
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 12986 7052 13806
rect 7208 13002 7236 20198
rect 7380 19780 7432 19786
rect 7380 19722 7432 19728
rect 7392 19174 7420 19722
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7484 18834 7512 20266
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7576 18426 7604 20470
rect 8024 20460 8076 20466
rect 8128 20448 8156 22200
rect 8076 20420 8156 20448
rect 8208 20460 8260 20466
rect 8024 20402 8076 20408
rect 8312 20448 8340 22222
rect 8588 22114 8616 22222
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 11978 22200 12034 23000
rect 12530 22200 12586 23000
rect 13082 22200 13138 23000
rect 13634 22200 13690 23000
rect 14186 22200 14242 23000
rect 14738 22200 14794 23000
rect 15290 22200 15346 23000
rect 15842 22200 15898 23000
rect 16394 22200 16450 23000
rect 16946 22200 17002 23000
rect 17498 22200 17554 23000
rect 18050 22200 18106 23000
rect 18602 22200 18658 23000
rect 19154 22200 19210 23000
rect 19706 22200 19762 23000
rect 20258 22200 20314 23000
rect 20810 22200 20866 23000
rect 21362 22200 21418 23000
rect 21560 22222 21864 22250
rect 8680 22114 8708 22200
rect 8588 22086 8708 22114
rect 9232 20534 9260 22200
rect 9784 20584 9812 22200
rect 9600 20556 9812 20584
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 8260 20420 8340 20448
rect 8208 20402 8260 20408
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7470 16552 7526 16561
rect 7470 16487 7526 16496
rect 7484 16454 7512 16487
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7300 16250 7328 16390
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7668 15570 7696 20198
rect 7760 17746 7788 20198
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7944 19514 7972 19654
rect 8036 19514 8064 19858
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8220 19446 8248 20402
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 9140 20058 9168 20266
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 8852 19984 8904 19990
rect 9036 19984 9088 19990
rect 8904 19932 9036 19938
rect 8852 19926 9088 19932
rect 8864 19910 9076 19926
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7852 16522 7880 18566
rect 8220 18290 8248 19246
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13530 7420 14214
rect 7576 14074 7604 14350
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7208 12986 7328 13002
rect 7012 12980 7064 12986
rect 7208 12980 7340 12986
rect 7208 12974 7288 12980
rect 7012 12922 7064 12928
rect 7288 12922 7340 12928
rect 7852 9450 7880 16458
rect 7944 15094 7972 16594
rect 8036 16454 8064 17002
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 8312 14074 8340 19314
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8404 17338 8432 18090
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8404 16250 8432 16390
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8496 16153 8524 19654
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17542 8616 18022
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8482 16144 8538 16153
rect 8482 16079 8538 16088
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8036 12102 8064 12786
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 10674 8064 12038
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10470 8064 10610
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7852 8838 7880 9386
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 8036 8362 8064 10406
rect 8128 8974 8156 13874
rect 8404 13258 8432 15302
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 12238 8248 12718
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11762 8248 12038
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8312 11642 8340 12174
rect 8680 11898 8708 19790
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9232 18970 9260 20470
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9324 18737 9352 20198
rect 9416 20058 9444 20334
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9508 19938 9536 20402
rect 9416 19910 9536 19938
rect 9416 18902 9444 19910
rect 9600 19854 9628 20556
rect 10336 20466 10364 22200
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 9678 20360 9734 20369
rect 9678 20295 9680 20304
rect 9732 20295 9734 20304
rect 9680 20266 9732 20272
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9600 19514 9628 19790
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9310 18728 9366 18737
rect 9310 18663 9366 18672
rect 9416 18630 9444 18838
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9140 15910 9168 17682
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8220 11614 8340 11642
rect 8220 10606 8248 11614
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8220 9042 8248 10542
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8312 9722 8340 10474
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 9178 8616 9522
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9140 6730 9168 15846
rect 9416 9586 9444 18566
rect 9692 18290 9720 19314
rect 9784 19242 9812 20402
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9876 19378 9904 19926
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17882 9812 18022
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16726 9812 16934
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9784 15502 9812 16526
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9600 14074 9628 15030
rect 9784 15026 9812 15438
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 10060 13530 10088 15370
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 12646 9812 13194
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 10152 12306 10180 12786
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 10674 9812 12038
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 9178 9444 9522
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9416 8838 9444 9114
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9968 6186 9996 9930
rect 10428 9654 10456 20538
rect 10888 20466 10916 22200
rect 11440 20890 11468 22200
rect 11256 20862 11468 20890
rect 11256 20466 11284 20862
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11992 20602 12020 22200
rect 12544 20602 12572 22200
rect 13096 20602 13124 22200
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10520 18426 10548 20198
rect 10704 18970 10732 20402
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10980 18698 11008 19790
rect 11072 18970 11100 20402
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19378 11192 19654
rect 11256 19446 11284 19790
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11716 19514 11744 19722
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10428 8906 10456 9590
rect 10520 9178 10548 12106
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10704 9042 10732 9318
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10796 8922 10824 18022
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10888 16046 10916 17138
rect 11256 16454 11284 18634
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11808 18358 11836 19450
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11900 19174 11928 19382
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18630 11928 19110
rect 12084 18630 12112 19178
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11900 18290 11928 18566
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11900 18086 11928 18226
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11900 16998 11928 18022
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16590 11928 16934
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 14890 10916 15982
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 11072 14482 11100 15302
rect 11256 14822 11284 16390
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15502 11560 15846
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11716 14890 11744 16458
rect 11900 16046 11928 16526
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11900 15910 11928 15982
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 14006 11100 14418
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14074 11284 14214
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11624 13530 11652 14010
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11624 13274 11652 13466
rect 11624 13246 11744 13274
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11716 12986 11744 13246
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11716 12102 11744 12922
rect 11808 12646 11836 13942
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11716 11150 11744 12038
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 9518 10916 10610
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10704 8894 10824 8922
rect 10888 8922 10916 9454
rect 10980 9110 11008 10406
rect 11900 10198 11928 13194
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11992 12986 12020 13126
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12084 12442 12112 13126
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11900 9110 11928 10134
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 10888 8894 11008 8922
rect 10704 8430 10732 8894
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8634 10824 8774
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10980 8430 11008 8894
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11164 8634 11192 8774
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10888 8242 10916 8366
rect 10888 8214 11100 8242
rect 11072 8022 11100 8214
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11256 7954 11284 8434
rect 11716 8090 11744 8502
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11808 5137 11836 8774
rect 12084 8022 12112 8842
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11900 6322 11928 7414
rect 12176 6914 12204 20198
rect 12452 19786 12480 20198
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12544 19174 12572 20402
rect 12728 19922 12756 20402
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12636 19446 12664 19790
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 13004 19378 13032 20334
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 13096 19922 13124 20266
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19922 13492 20198
rect 13556 20058 13584 20334
rect 13648 20074 13676 22200
rect 14200 20330 14228 22200
rect 14752 20602 14780 22200
rect 14740 20596 14792 20602
rect 15304 20584 15332 22200
rect 15384 20596 15436 20602
rect 15304 20556 15384 20584
rect 14740 20538 14792 20544
rect 15856 20584 15884 22200
rect 15936 20596 15988 20602
rect 15856 20556 15936 20584
rect 15384 20538 15436 20544
rect 15936 20538 15988 20544
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 13648 20058 13860 20074
rect 14660 20058 14688 20402
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 13544 20052 13596 20058
rect 13648 20052 13872 20058
rect 13648 20046 13820 20052
rect 13544 19994 13596 20000
rect 13820 19994 13872 20000
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 15304 19990 15332 20334
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14832 19848 14884 19854
rect 15108 19848 15160 19854
rect 14832 19790 14884 19796
rect 15106 19816 15108 19825
rect 15160 19816 15162 19825
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12268 16250 12296 16458
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12268 15026 12296 15642
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 15094 12388 15438
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12360 10742 12388 11086
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12360 10266 12388 10678
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8634 12296 8774
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12452 8430 12480 11086
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12176 6886 12388 6914
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12360 6118 12388 6886
rect 12544 6225 12572 19110
rect 12728 18358 12756 19314
rect 13188 18630 13216 19654
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13004 16182 13032 16934
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12820 14074 12848 15370
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12820 13802 12848 14010
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 13556 12434 13584 18566
rect 13832 17202 13860 18702
rect 14384 18086 14412 19110
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14292 17270 14320 18022
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 16454 13860 17138
rect 14384 17134 14412 18022
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14384 16658 14412 17070
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 14384 16250 14412 16594
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 14292 13870 14320 14758
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13832 12646 13860 12922
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13464 12406 13584 12434
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 6254 12940 10542
rect 13004 10470 13032 11018
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12900 6248 12952 6254
rect 12530 6216 12586 6225
rect 12900 6190 12952 6196
rect 12530 6151 12586 6160
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12912 5778 12940 6190
rect 13004 6186 13032 10406
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8634 13216 8774
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 13464 5166 13492 12406
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 11898 13952 12174
rect 14292 12102 14320 12786
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10674 13768 10950
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13832 9994 13860 11290
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 8838 13584 9522
rect 13832 9042 13860 9930
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8634 13584 8774
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 6866 13676 7142
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6186 13768 6734
rect 13832 6662 13860 7822
rect 14292 7274 14320 12038
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 6390 13952 6598
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14384 6254 14412 10406
rect 14476 10062 14504 19790
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 14006 14688 14214
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14844 13258 14872 19790
rect 15106 19751 15162 19760
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15304 15910 15332 16118
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13326 15056 13670
rect 15304 13326 15332 15846
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 15028 12918 15056 13262
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12434 14964 12582
rect 14844 12406 14964 12434
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14568 11354 14596 12242
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8566 14504 8774
rect 14660 8634 14688 9386
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14660 7750 14688 8570
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14660 6186 14688 6802
rect 14844 6730 14872 12406
rect 15028 12238 15056 12854
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10470 15056 10950
rect 15120 10742 15148 11018
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15120 10606 15148 10678
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15120 10266 15148 10542
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9042 15424 9318
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 8634 14964 8774
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15212 7886 15240 8298
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14936 6866 14964 7210
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14844 6458 14872 6666
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14660 5234 14688 6122
rect 14844 6100 14872 6394
rect 14924 6112 14976 6118
rect 14844 6072 14924 6100
rect 14924 6054 14976 6060
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 13452 5160 13504 5166
rect 11794 5128 11850 5137
rect 13452 5102 13504 5108
rect 11794 5063 11850 5072
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 15028 2854 15056 7686
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6662 15240 7142
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5914 15148 6258
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15212 4282 15240 6326
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 15212 2514 15240 4218
rect 15304 3670 15332 8502
rect 15396 4826 15424 8978
rect 15488 8430 15516 20402
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 17202 15884 19654
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15948 17678 15976 18158
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 16040 17338 16068 19382
rect 16132 17882 16160 19790
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15856 14346 15884 15302
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15580 5370 15608 5510
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15672 5302 15700 6598
rect 15764 6458 15792 6598
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15856 4078 15884 14282
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16132 10266 16160 12106
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16132 8974 16160 10202
rect 16224 9382 16252 20402
rect 16408 20244 16436 22200
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16960 20330 16988 22200
rect 17512 20602 17540 22200
rect 17500 20596 17552 20602
rect 18064 20584 18092 22200
rect 18064 20556 18184 20584
rect 17500 20538 17552 20544
rect 17958 20496 18014 20505
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17592 20460 17644 20466
rect 17958 20431 18014 20440
rect 18052 20460 18104 20466
rect 17592 20402 17644 20408
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16580 20256 16632 20262
rect 16408 20216 16580 20244
rect 16580 20198 16632 20204
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16408 17882 16436 19722
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16868 17814 16896 18294
rect 16960 18290 16988 18566
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16960 17338 16988 18226
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 17052 16232 17080 20402
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 16960 16204 17080 16232
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16408 13530 16436 15370
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16684 14618 16712 14962
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16408 13274 16436 13466
rect 16316 13246 16436 13274
rect 16316 12866 16344 13246
rect 16488 13184 16540 13190
rect 16408 13144 16488 13172
rect 16408 12986 16436 13144
rect 16488 13126 16540 13132
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16316 12838 16436 12866
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8498 16252 8774
rect 16316 8634 16344 8842
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 6458 15976 7142
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16408 4622 16436 12838
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16684 9994 16712 10542
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 7993 16988 16204
rect 17144 15162 17172 19790
rect 17236 19514 17264 19858
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18358 17264 19110
rect 17420 18766 17448 19654
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17512 17542 17540 17818
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17512 14618 17540 14962
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17052 13462 17080 14282
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12646 17080 13194
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16946 7984 17002 7993
rect 16946 7919 17002 7928
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 17052 6866 17080 12582
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8634 17172 8910
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17420 6662 17448 8366
rect 17512 8090 17540 8434
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 17236 6474 17264 6598
rect 17236 6446 17356 6474
rect 17512 6458 17540 6666
rect 17328 6390 17356 6446
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17604 5846 17632 20402
rect 17972 20210 18000 20431
rect 18052 20402 18104 20408
rect 17788 20182 18000 20210
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17696 17066 17724 19790
rect 17788 19718 17816 20182
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17880 19378 17908 19994
rect 18064 19417 18092 20402
rect 18156 20330 18184 20556
rect 18418 20360 18474 20369
rect 18144 20324 18196 20330
rect 18418 20295 18474 20304
rect 18144 20266 18196 20272
rect 18432 19922 18460 20295
rect 18616 20058 18644 22200
rect 18970 21040 19026 21049
rect 18970 20975 19026 20984
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18510 19952 18566 19961
rect 18420 19916 18472 19922
rect 18510 19887 18566 19896
rect 18604 19916 18656 19922
rect 18420 19858 18472 19864
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18050 19408 18106 19417
rect 17868 19372 17920 19378
rect 18050 19343 18106 19352
rect 17868 19314 17920 19320
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18086 17908 18566
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17880 17746 17908 18022
rect 17972 17882 18000 19178
rect 18064 18970 18092 19246
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18248 18766 18276 19654
rect 18524 19378 18552 19887
rect 18604 19858 18656 19864
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 18616 17610 18644 19858
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18892 18902 18920 19314
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 18616 16794 18644 17546
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18144 16584 18196 16590
rect 17958 16552 18014 16561
rect 18144 16526 18196 16532
rect 17958 16487 18014 16496
rect 17972 16114 18000 16487
rect 18156 16153 18184 16526
rect 18142 16144 18198 16153
rect 17960 16108 18012 16114
rect 18142 16079 18198 16088
rect 17960 16050 18012 16056
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 17696 15570 17724 15846
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 18248 15502 18276 15846
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 14414 17908 15302
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 13870 17908 14350
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 13530 17908 13806
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17880 7954 17908 10474
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17880 7834 17908 7890
rect 17788 7806 17908 7834
rect 17788 6866 17816 7806
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17696 6458 17724 6598
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17880 5914 17908 7686
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 4146 16436 4558
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 17052 4282 17080 4422
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 17972 2922 18000 8298
rect 18064 6662 18092 13194
rect 18708 13190 18736 18770
rect 18984 18426 19012 20975
rect 19168 20584 19196 22200
rect 19340 20596 19392 20602
rect 19168 20556 19340 20584
rect 19340 20538 19392 20544
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19062 19816 19118 19825
rect 19062 19751 19118 19760
rect 19076 19378 19104 19751
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19156 19304 19208 19310
rect 19076 19252 19156 19258
rect 19076 19246 19208 19252
rect 19076 19230 19196 19246
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18800 16114 18828 16662
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18800 12850 18828 14214
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18156 8634 18184 9590
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18248 6254 18276 10746
rect 18340 10470 18368 11018
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 8430 18368 10406
rect 18418 9752 18474 9761
rect 18418 9687 18474 9696
rect 18432 9654 18460 9687
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18156 6118 18184 6190
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5914 18184 6054
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18248 5778 18276 6190
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18248 5030 18276 5510
rect 18340 5302 18368 5578
rect 18708 5545 18736 11834
rect 18800 11642 18828 12786
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 11778 18920 12582
rect 18984 11898 19012 18226
rect 19076 15706 19104 19230
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19536 18290 19564 20266
rect 19628 19666 19656 20470
rect 19720 20330 19748 22200
rect 20272 20602 20300 22200
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19708 20324 19760 20330
rect 19708 20266 19760 20272
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19628 19638 19748 19666
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19628 19417 19656 19450
rect 19614 19408 19670 19417
rect 19614 19343 19670 19352
rect 19720 18442 19748 19638
rect 19812 18834 19840 19858
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19628 18414 19748 18442
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19352 17338 19380 17682
rect 19628 17626 19656 18414
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19536 17598 19656 17626
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19536 17082 19564 17598
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19628 17202 19656 17478
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19536 17054 19656 17082
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19536 16454 19564 16934
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19536 13938 19564 14554
rect 19628 14278 19656 17054
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19536 13530 19564 13874
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19536 12986 19564 13466
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18892 11750 19012 11778
rect 18800 11614 18920 11642
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11150 18828 11494
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18892 8362 18920 11614
rect 18984 11098 19012 11750
rect 19076 11257 19104 12038
rect 19536 11558 19564 12922
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19062 11248 19118 11257
rect 19062 11183 19118 11192
rect 18984 11082 19104 11098
rect 18984 11076 19116 11082
rect 18984 11070 19064 11076
rect 19064 11018 19116 11024
rect 19076 9042 19104 11018
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19246 9072 19302 9081
rect 19064 9036 19116 9042
rect 19246 9007 19302 9016
rect 19064 8978 19116 8984
rect 19260 8974 19288 9007
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 19076 8294 19104 8774
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19260 7546 19288 7890
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19536 6458 19564 10066
rect 19628 6866 19656 11494
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18694 5536 18750 5545
rect 18694 5471 18750 5480
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4078 18276 4966
rect 18340 4758 18368 5238
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 18340 4486 18368 4694
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 18800 2774 18828 5850
rect 18892 5817 18920 6258
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 18878 5808 18934 5817
rect 19076 5778 19104 6054
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19246 5808 19302 5817
rect 18878 5743 18934 5752
rect 19064 5772 19116 5778
rect 19246 5743 19302 5752
rect 19064 5714 19116 5720
rect 19260 5370 19288 5743
rect 19536 5574 19564 6122
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4010 19288 4558
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19536 3194 19564 5510
rect 19720 4826 19748 18226
rect 19812 18154 19840 18770
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19812 17678 19840 18090
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19812 14822 19840 16050
rect 19904 15706 19932 20402
rect 20824 19530 20852 22200
rect 21086 21448 21142 21457
rect 21086 21383 21142 21392
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20640 19514 20852 19530
rect 20628 19508 20852 19514
rect 20680 19502 20852 19508
rect 20628 19450 20680 19456
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19904 11558 19932 13942
rect 19996 12986 20024 19314
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 19009 20760 19110
rect 20718 19000 20774 19009
rect 20718 18935 20774 18944
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20166 18184 20222 18193
rect 20166 18119 20168 18128
rect 20220 18119 20222 18128
rect 20168 18090 20220 18096
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20088 16250 20116 17138
rect 20168 16992 20220 16998
rect 20166 16960 20168 16969
rect 20220 16960 20222 16969
rect 20166 16895 20222 16904
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19812 10674 19840 11018
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19812 9994 19840 10610
rect 20088 10266 20116 14350
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 9988 19852 9994
rect 19800 9930 19852 9936
rect 19904 9625 19932 9998
rect 19890 9616 19946 9625
rect 19800 9580 19852 9586
rect 19890 9551 19946 9560
rect 19800 9522 19852 9528
rect 19812 9217 19840 9522
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19798 9208 19854 9217
rect 19798 9143 19854 9152
rect 19812 9042 19840 9143
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 5914 19840 8434
rect 19904 7818 19932 8570
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19904 6390 19932 7754
rect 19996 6866 20024 9386
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 20088 7546 20116 8774
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20180 7274 20208 15098
rect 20272 13530 20300 18634
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20364 14226 20392 15982
rect 20456 15706 20484 18226
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17785 20668 18022
rect 20626 17776 20682 17785
rect 20626 17711 20682 17720
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 16561 20576 16934
rect 20640 16794 20668 17546
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20534 16552 20590 16561
rect 20534 16487 20590 16496
rect 20640 16250 20668 16730
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20548 15162 20576 16050
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20640 14618 20668 16186
rect 20732 16182 20760 17138
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15745 20760 15846
rect 20718 15736 20774 15745
rect 20718 15671 20774 15680
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20364 14198 20484 14226
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 12889 20392 13262
rect 20350 12880 20406 12889
rect 20260 12844 20312 12850
rect 20350 12815 20406 12824
rect 20260 12786 20312 12792
rect 20272 12442 20300 12786
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20350 10432 20406 10441
rect 20350 10367 20406 10376
rect 20364 10062 20392 10367
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20364 9722 20392 9998
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 9178 20300 9522
rect 20456 9450 20484 14198
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20548 12374 20576 12786
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20444 9444 20496 9450
rect 20444 9386 20496 9392
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20548 8974 20576 9862
rect 20640 9042 20668 13874
rect 20732 9450 20760 15370
rect 20824 14890 20852 19314
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20824 11914 20852 14010
rect 20916 12442 20944 20402
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21008 13410 21036 20334
rect 21100 19854 21128 21383
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 21086 18728 21142 18737
rect 21086 18663 21142 18672
rect 21100 18630 21128 18663
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21100 17338 21128 18226
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21192 14074 21220 20470
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18737 21312 19110
rect 21376 18970 21404 22200
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21270 18728 21326 18737
rect 21560 18698 21588 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22466 22200 22522 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21270 18663 21326 18672
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21284 17241 21312 18022
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21284 16153 21312 16934
rect 21376 16590 21404 18566
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 22480 18154 22508 22200
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21270 16144 21326 16153
rect 21270 16079 21326 16088
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15473 21312 15846
rect 22192 15496 22244 15502
rect 21270 15464 21326 15473
rect 22192 15438 22244 15444
rect 21270 15399 21326 15408
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21284 14929 21312 15302
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21270 14920 21326 14929
rect 21270 14855 21326 14864
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21284 14521 21312 14758
rect 21270 14512 21326 14521
rect 21270 14447 21326 14456
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21284 13977 21312 14214
rect 21270 13968 21326 13977
rect 21270 13903 21326 13912
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21270 13696 21326 13705
rect 21270 13631 21326 13640
rect 21284 13530 21312 13631
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21008 13382 21128 13410
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21008 12442 21036 13262
rect 21100 12986 21128 13382
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21270 13288 21326 13297
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20824 11886 20944 11914
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20824 11286 20852 11766
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20548 8634 20576 8774
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20364 8401 20392 8434
rect 20350 8392 20406 8401
rect 20350 8327 20406 8336
rect 20364 8090 20392 8327
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20732 8106 20760 8230
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20548 8078 20760 8106
rect 20548 8022 20576 8078
rect 20536 8016 20588 8022
rect 20720 8016 20772 8022
rect 20536 7958 20588 7964
rect 20718 7984 20720 7993
rect 20772 7984 20774 7993
rect 20718 7919 20774 7928
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20350 7168 20406 7177
rect 20350 7103 20406 7112
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 20364 6798 20392 7103
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20718 6760 20774 6769
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6458 20300 6598
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 19892 6384 19944 6390
rect 19892 6326 19944 6332
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19996 5710 20024 6287
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19996 5370 20024 5646
rect 20364 5370 20392 6734
rect 20718 6695 20774 6704
rect 20732 6662 20760 6695
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20640 6458 20668 6598
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20548 5914 20576 6326
rect 20824 6254 20852 11222
rect 20916 10810 20944 11886
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20902 10024 20958 10033
rect 20902 9959 20958 9968
rect 20916 9586 20944 9959
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21008 8616 21036 9454
rect 21100 9178 21128 12786
rect 21192 12434 21220 13262
rect 21270 13223 21326 13232
rect 21284 12986 21312 13223
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21376 12481 21404 12582
rect 21362 12472 21418 12481
rect 21192 12406 21312 12434
rect 21362 12407 21418 12416
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21192 11354 21220 12174
rect 21284 11830 21312 12406
rect 21376 12238 21404 12407
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21272 11688 21324 11694
rect 21376 11665 21404 11698
rect 21272 11630 21324 11636
rect 21362 11656 21418 11665
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21284 10742 21312 11630
rect 21362 11591 21418 11600
rect 21376 11150 21404 11591
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 10736 21324 10742
rect 21178 10704 21234 10713
rect 21272 10678 21324 10684
rect 21178 10639 21234 10648
rect 21192 9761 21220 10639
rect 21284 9926 21312 10678
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21178 9752 21234 9761
rect 21178 9687 21234 9696
rect 21192 9586 21220 9687
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21284 8634 21312 9862
rect 21468 9450 21496 13874
rect 21546 12200 21602 12209
rect 21546 12135 21548 12144
rect 21600 12135 21602 12144
rect 21548 12106 21600 12112
rect 21560 11898 21588 12106
rect 21652 12102 21680 14350
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21362 8936 21418 8945
rect 21362 8871 21418 8880
rect 21272 8628 21324 8634
rect 21008 8588 21128 8616
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20916 7886 20944 8298
rect 21008 8090 21036 8434
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21008 7750 21036 7822
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21100 7546 21128 8588
rect 21272 8570 21324 8576
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21192 7886 21220 7958
rect 21376 7886 21404 8871
rect 21454 7984 21510 7993
rect 21454 7919 21510 7928
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20812 6248 20864 6254
rect 20718 6216 20774 6225
rect 20812 6190 20864 6196
rect 20718 6151 20774 6160
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20732 5846 20760 6151
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20442 5536 20498 5545
rect 20442 5471 20498 5480
rect 20626 5536 20682 5545
rect 20626 5471 20682 5480
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20350 5128 20406 5137
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 20088 4690 20116 4966
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20272 4282 20300 5102
rect 20350 5063 20352 5072
rect 20404 5063 20406 5072
rect 20352 5034 20404 5040
rect 20456 4826 20484 5471
rect 20640 5302 20668 5471
rect 20628 5296 20680 5302
rect 20548 5244 20628 5250
rect 20548 5238 20680 5244
rect 20548 5222 20668 5238
rect 20824 5234 20852 6054
rect 21192 5642 21220 7686
rect 21376 7449 21404 7686
rect 21362 7440 21418 7449
rect 21468 7410 21496 7919
rect 21362 7375 21418 7384
rect 21456 7404 21508 7410
rect 21376 6866 21404 7375
rect 21456 7346 21508 7352
rect 21560 7342 21588 10542
rect 21652 8294 21680 11766
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 22112 8906 22140 14962
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21362 6760 21418 6769
rect 21362 6695 21418 6704
rect 21376 6458 21404 6695
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 20812 5228 20864 5234
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20350 4720 20406 4729
rect 20350 4655 20406 4664
rect 20364 4622 20392 4655
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20166 3904 20222 3913
rect 20166 3839 20222 3848
rect 20180 3738 20208 3839
rect 20364 3738 20392 4558
rect 20548 4282 20576 5222
rect 20812 5170 20864 5176
rect 20628 5160 20680 5166
rect 20626 5128 20628 5137
rect 20680 5128 20682 5137
rect 22204 5098 22232 15438
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22296 8022 22324 12038
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 20626 5063 20682 5072
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21376 4282 21404 4490
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21272 4208 21324 4214
rect 21376 4185 21404 4218
rect 21272 4150 21324 4156
rect 21362 4176 21418 4185
rect 21284 3913 21312 4150
rect 21362 4111 21418 4120
rect 21270 3904 21326 3913
rect 21270 3839 21326 3848
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 21270 3496 21326 3505
rect 21270 3431 21272 3440
rect 21324 3431 21326 3440
rect 21272 3402 21324 3408
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 21270 3088 21326 3097
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 18800 2746 18920 2774
rect 18892 2582 18920 2746
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 20166 2408 20222 2417
rect 20166 2343 20168 2352
rect 20220 2343 20222 2352
rect 20168 2314 20220 2320
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 20272 1873 20300 2994
rect 20640 2689 20668 3062
rect 21270 3023 21272 3032
rect 21324 3023 21326 3032
rect 21272 2994 21324 3000
rect 20626 2680 20682 2689
rect 20626 2615 20682 2624
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20258 1864 20314 1873
rect 20258 1799 20314 1808
rect 20548 1465 20576 2382
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 20534 1456 20590 1465
rect 20534 1391 20590 1400
<< via2 >>
rect 1490 17176 1546 17232
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5446 9016 5502 9072
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 1398 5752 1454 5808
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6918 19760 6974 19816
rect 7470 16496 7526 16552
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8482 16088 8538 16144
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 9678 20324 9734 20360
rect 9678 20304 9680 20324
rect 9680 20304 9732 20324
rect 9732 20304 9734 20324
rect 9310 18672 9366 18728
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 15106 19796 15108 19816
rect 15108 19796 15160 19816
rect 15160 19796 15162 19816
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 12530 6160 12586 6216
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 15106 19760 15162 19796
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 11794 5072 11850 5128
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 17958 20440 18014 20496
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16946 7928 17002 7984
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 18418 20304 18474 20360
rect 18970 20984 19026 21040
rect 18510 19896 18566 19952
rect 18050 19352 18106 19408
rect 17958 16496 18014 16552
rect 18142 16088 18198 16144
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19062 19760 19118 19816
rect 18418 9696 18474 9752
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19614 19352 19670 19408
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19062 11192 19118 11248
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19246 9016 19302 9072
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18694 5480 18750 5536
rect 18878 5752 18934 5808
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19246 5752 19302 5808
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 21086 21392 21142 21448
rect 20718 18944 20774 19000
rect 20166 18148 20222 18184
rect 20166 18128 20168 18148
rect 20168 18128 20220 18148
rect 20220 18128 20222 18148
rect 20166 16940 20168 16960
rect 20168 16940 20220 16960
rect 20220 16940 20222 16960
rect 20166 16904 20222 16940
rect 19890 9560 19946 9616
rect 19798 9152 19854 9208
rect 20626 17720 20682 17776
rect 20534 16496 20590 16552
rect 20718 15680 20774 15736
rect 20350 12824 20406 12880
rect 20350 10376 20406 10432
rect 21086 18672 21142 18728
rect 21270 18672 21326 18728
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21270 17176 21326 17232
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21270 16088 21326 16144
rect 21270 15408 21326 15464
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21270 14864 21326 14920
rect 21270 14456 21326 14512
rect 21270 13912 21326 13968
rect 21270 13640 21326 13696
rect 20350 8336 20406 8392
rect 20718 7964 20720 7984
rect 20720 7964 20772 7984
rect 20772 7964 20774 7984
rect 20718 7928 20774 7964
rect 20350 7112 20406 7168
rect 19982 6296 20038 6352
rect 20718 6704 20774 6760
rect 20902 9968 20958 10024
rect 21270 13232 21326 13288
rect 21362 12416 21418 12472
rect 21362 11600 21418 11656
rect 21178 10648 21234 10704
rect 21178 9696 21234 9752
rect 21546 12164 21602 12200
rect 21546 12144 21548 12164
rect 21548 12144 21600 12164
rect 21600 12144 21602 12164
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21362 8880 21418 8936
rect 21454 7928 21510 7984
rect 20718 6160 20774 6216
rect 20442 5480 20498 5536
rect 20626 5480 20682 5536
rect 20350 5092 20406 5128
rect 20350 5072 20352 5092
rect 20352 5072 20404 5092
rect 20404 5072 20406 5092
rect 21362 7384 21418 7440
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21362 6704 21418 6760
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 20350 4664 20406 4720
rect 20166 3848 20222 3904
rect 20626 5108 20628 5128
rect 20628 5108 20680 5128
rect 20680 5108 20682 5128
rect 20626 5072 20682 5108
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21362 4120 21418 4176
rect 21270 3848 21326 3904
rect 21270 3460 21326 3496
rect 21270 3440 21272 3460
rect 21272 3440 21324 3460
rect 21324 3440 21326 3460
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 20166 2372 20222 2408
rect 20166 2352 20168 2372
rect 20168 2352 20220 2372
rect 20220 2352 20222 2372
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 21270 3052 21326 3088
rect 21270 3032 21272 3052
rect 21272 3032 21324 3052
rect 21324 3032 21326 3052
rect 20626 2624 20682 2680
rect 20258 1808 20314 1864
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 20534 1400 20590 1456
<< metal3 >>
rect 21081 21450 21147 21453
rect 22200 21450 23000 21480
rect 21081 21448 23000 21450
rect 21081 21392 21086 21448
rect 21142 21392 23000 21448
rect 21081 21390 23000 21392
rect 21081 21387 21147 21390
rect 22200 21360 23000 21390
rect 18965 21042 19031 21045
rect 22200 21042 23000 21072
rect 18965 21040 23000 21042
rect 18965 20984 18970 21040
rect 19026 20984 23000 21040
rect 18965 20982 23000 20984
rect 18965 20979 19031 20982
rect 22200 20952 23000 20982
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 22200 20634 23000 20664
rect 22142 20544 23000 20634
rect 17953 20498 18019 20501
rect 22142 20498 22202 20544
rect 17953 20496 22202 20498
rect 17953 20440 17958 20496
rect 18014 20440 22202 20496
rect 17953 20438 22202 20440
rect 17953 20435 18019 20438
rect 9673 20362 9739 20365
rect 18413 20362 18479 20365
rect 9673 20360 18479 20362
rect 9673 20304 9678 20360
rect 9734 20304 18418 20360
rect 18474 20304 18479 20360
rect 9673 20302 18479 20304
rect 9673 20299 9739 20302
rect 18413 20299 18479 20302
rect 22200 20226 23000 20256
rect 19934 20166 23000 20226
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 18505 19954 18571 19957
rect 19934 19954 19994 20166
rect 22200 20136 23000 20166
rect 18505 19952 19994 19954
rect 18505 19896 18510 19952
rect 18566 19896 19994 19952
rect 18505 19894 19994 19896
rect 18505 19891 18571 19894
rect 6913 19818 6979 19821
rect 15101 19818 15167 19821
rect 6913 19816 15167 19818
rect 6913 19760 6918 19816
rect 6974 19760 15106 19816
rect 15162 19760 15167 19816
rect 6913 19758 15167 19760
rect 6913 19755 6979 19758
rect 15101 19755 15167 19758
rect 19057 19818 19123 19821
rect 22200 19818 23000 19848
rect 19057 19816 23000 19818
rect 19057 19760 19062 19816
rect 19118 19760 23000 19816
rect 19057 19758 23000 19760
rect 19057 19755 19123 19758
rect 22200 19728 23000 19758
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 18045 19412 18111 19413
rect 18045 19408 18092 19412
rect 18156 19410 18162 19412
rect 19609 19410 19675 19413
rect 22200 19410 23000 19440
rect 18045 19352 18050 19408
rect 18045 19348 18092 19352
rect 18156 19350 18202 19410
rect 19609 19408 23000 19410
rect 19609 19352 19614 19408
rect 19670 19352 23000 19408
rect 19609 19350 23000 19352
rect 18156 19348 18162 19350
rect 18045 19347 18111 19348
rect 19609 19347 19675 19350
rect 22200 19320 23000 19350
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 20713 19002 20779 19005
rect 22200 19002 23000 19032
rect 20713 19000 23000 19002
rect 20713 18944 20718 19000
rect 20774 18944 23000 19000
rect 20713 18942 23000 18944
rect 20713 18939 20779 18942
rect 22200 18912 23000 18942
rect 9305 18730 9371 18733
rect 21081 18730 21147 18733
rect 9305 18728 21147 18730
rect 9305 18672 9310 18728
rect 9366 18672 21086 18728
rect 21142 18672 21147 18728
rect 9305 18670 21147 18672
rect 9305 18667 9371 18670
rect 21081 18667 21147 18670
rect 21265 18730 21331 18733
rect 21265 18728 22202 18730
rect 21265 18672 21270 18728
rect 21326 18672 22202 18728
rect 21265 18670 22202 18672
rect 21265 18667 21331 18670
rect 22142 18624 22202 18670
rect 22142 18534 23000 18624
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 20161 18186 20227 18189
rect 22200 18186 23000 18216
rect 20161 18184 23000 18186
rect 20161 18128 20166 18184
rect 20222 18128 23000 18184
rect 20161 18126 23000 18128
rect 20161 18123 20227 18126
rect 22200 18096 23000 18126
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 20621 17778 20687 17781
rect 22200 17778 23000 17808
rect 20621 17776 23000 17778
rect 20621 17720 20626 17776
rect 20682 17720 23000 17776
rect 20621 17718 23000 17720
rect 20621 17715 20687 17718
rect 22200 17688 23000 17718
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 22200 17370 23000 17400
rect 22142 17280 23000 17370
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 21265 17234 21331 17237
rect 22142 17234 22202 17280
rect 21265 17232 22202 17234
rect 21265 17176 21270 17232
rect 21326 17176 22202 17232
rect 21265 17174 22202 17176
rect 21265 17171 21331 17174
rect 20161 16962 20227 16965
rect 22200 16962 23000 16992
rect 20161 16960 23000 16962
rect 20161 16904 20166 16960
rect 20222 16904 23000 16960
rect 20161 16902 23000 16904
rect 20161 16899 20227 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 7465 16554 7531 16557
rect 17953 16554 18019 16557
rect 7465 16552 18019 16554
rect 7465 16496 7470 16552
rect 7526 16496 17958 16552
rect 18014 16496 18019 16552
rect 7465 16494 18019 16496
rect 7465 16491 7531 16494
rect 17953 16491 18019 16494
rect 20529 16554 20595 16557
rect 22200 16554 23000 16584
rect 20529 16552 23000 16554
rect 20529 16496 20534 16552
rect 20590 16496 23000 16552
rect 20529 16494 23000 16496
rect 20529 16491 20595 16494
rect 22200 16464 23000 16494
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 8477 16146 8543 16149
rect 18137 16146 18203 16149
rect 8477 16144 18203 16146
rect 8477 16088 8482 16144
rect 8538 16088 18142 16144
rect 18198 16088 18203 16144
rect 8477 16086 18203 16088
rect 8477 16083 8543 16086
rect 18137 16083 18203 16086
rect 21265 16146 21331 16149
rect 22200 16146 23000 16176
rect 21265 16144 23000 16146
rect 21265 16088 21270 16144
rect 21326 16088 23000 16144
rect 21265 16086 23000 16088
rect 21265 16083 21331 16086
rect 22200 16056 23000 16086
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 20713 15738 20779 15741
rect 22200 15738 23000 15768
rect 20713 15736 23000 15738
rect 20713 15680 20718 15736
rect 20774 15680 23000 15736
rect 20713 15678 23000 15680
rect 20713 15675 20779 15678
rect 22200 15648 23000 15678
rect 21265 15466 21331 15469
rect 21265 15464 22202 15466
rect 21265 15408 21270 15464
rect 21326 15408 22202 15464
rect 21265 15406 22202 15408
rect 21265 15403 21331 15406
rect 22142 15360 22202 15406
rect 22142 15270 23000 15360
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 21265 14922 21331 14925
rect 22200 14922 23000 14952
rect 21265 14920 23000 14922
rect 21265 14864 21270 14920
rect 21326 14864 23000 14920
rect 21265 14862 23000 14864
rect 21265 14859 21331 14862
rect 22200 14832 23000 14862
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 21265 14514 21331 14517
rect 22200 14514 23000 14544
rect 21265 14512 23000 14514
rect 21265 14456 21270 14512
rect 21326 14456 23000 14512
rect 21265 14454 23000 14456
rect 21265 14451 21331 14454
rect 22200 14424 23000 14454
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 22200 14106 23000 14136
rect 22142 14016 23000 14106
rect 21265 13970 21331 13973
rect 22142 13970 22202 14016
rect 21265 13968 22202 13970
rect 21265 13912 21270 13968
rect 21326 13912 22202 13968
rect 21265 13910 22202 13912
rect 21265 13907 21331 13910
rect 21265 13698 21331 13701
rect 22200 13698 23000 13728
rect 21265 13696 23000 13698
rect 21265 13640 21270 13696
rect 21326 13640 23000 13696
rect 21265 13638 23000 13640
rect 21265 13635 21331 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22200 13608 23000 13638
rect 19139 13567 19455 13568
rect 21265 13290 21331 13293
rect 22200 13290 23000 13320
rect 21265 13288 23000 13290
rect 21265 13232 21270 13288
rect 21326 13232 23000 13288
rect 21265 13230 23000 13232
rect 21265 13227 21331 13230
rect 22200 13200 23000 13230
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 20345 12882 20411 12885
rect 22200 12882 23000 12912
rect 20345 12880 23000 12882
rect 20345 12824 20350 12880
rect 20406 12824 23000 12880
rect 20345 12822 23000 12824
rect 20345 12819 20411 12822
rect 22200 12792 23000 12822
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 21357 12474 21423 12477
rect 22200 12474 23000 12504
rect 21357 12472 23000 12474
rect 21357 12416 21362 12472
rect 21418 12416 23000 12472
rect 21357 12414 23000 12416
rect 21357 12411 21423 12414
rect 22200 12384 23000 12414
rect 21541 12202 21607 12205
rect 21541 12200 22202 12202
rect 21541 12144 21546 12200
rect 21602 12144 22202 12200
rect 21541 12142 22202 12144
rect 21541 12139 21607 12142
rect 22142 12096 22202 12142
rect 22142 12006 23000 12096
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 21357 11658 21423 11661
rect 22200 11658 23000 11688
rect 21357 11656 23000 11658
rect 21357 11600 21362 11656
rect 21418 11600 23000 11656
rect 21357 11598 23000 11600
rect 21357 11595 21423 11598
rect 22200 11568 23000 11598
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 19057 11250 19123 11253
rect 22200 11250 23000 11280
rect 19057 11248 23000 11250
rect 19057 11192 19062 11248
rect 19118 11192 23000 11248
rect 19057 11190 23000 11192
rect 19057 11187 19123 11190
rect 22200 11160 23000 11190
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 22200 10842 23000 10872
rect 22142 10752 23000 10842
rect 21173 10706 21239 10709
rect 22142 10706 22202 10752
rect 21173 10704 22202 10706
rect 21173 10648 21178 10704
rect 21234 10648 22202 10704
rect 21173 10646 22202 10648
rect 21173 10643 21239 10646
rect 20345 10434 20411 10437
rect 22200 10434 23000 10464
rect 20345 10432 23000 10434
rect 20345 10376 20350 10432
rect 20406 10376 23000 10432
rect 20345 10374 23000 10376
rect 20345 10371 20411 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 22200 10344 23000 10374
rect 19139 10303 19455 10304
rect 20897 10026 20963 10029
rect 22200 10026 23000 10056
rect 20897 10024 23000 10026
rect 20897 9968 20902 10024
rect 20958 9968 23000 10024
rect 20897 9966 23000 9968
rect 20897 9963 20963 9966
rect 22200 9936 23000 9966
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 18413 9754 18479 9757
rect 21173 9754 21239 9757
rect 18413 9752 21239 9754
rect 18413 9696 18418 9752
rect 18474 9696 21178 9752
rect 21234 9696 21239 9752
rect 18413 9694 21239 9696
rect 18413 9691 18479 9694
rect 21173 9691 21239 9694
rect 19885 9618 19951 9621
rect 22200 9618 23000 9648
rect 19885 9616 23000 9618
rect 19885 9560 19890 9616
rect 19946 9560 23000 9616
rect 19885 9558 23000 9560
rect 19885 9555 19951 9558
rect 22200 9528 23000 9558
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 19793 9210 19859 9213
rect 22200 9210 23000 9240
rect 19793 9208 23000 9210
rect 19793 9152 19798 9208
rect 19854 9152 23000 9208
rect 19793 9150 23000 9152
rect 19793 9147 19859 9150
rect 22200 9120 23000 9150
rect 5441 9074 5507 9077
rect 19241 9074 19307 9077
rect 5441 9072 19307 9074
rect 5441 9016 5446 9072
rect 5502 9016 19246 9072
rect 19302 9016 19307 9072
rect 5441 9014 19307 9016
rect 5441 9011 5507 9014
rect 19241 9011 19307 9014
rect 21357 8938 21423 8941
rect 21357 8936 22202 8938
rect 21357 8880 21362 8936
rect 21418 8880 22202 8936
rect 21357 8878 22202 8880
rect 21357 8875 21423 8878
rect 22142 8832 22202 8878
rect 22142 8742 23000 8832
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 20345 8394 20411 8397
rect 22200 8394 23000 8424
rect 20345 8392 23000 8394
rect 20345 8336 20350 8392
rect 20406 8336 23000 8392
rect 20345 8334 23000 8336
rect 20345 8331 20411 8334
rect 22200 8304 23000 8334
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 16941 7986 17007 7989
rect 20713 7986 20779 7989
rect 16941 7984 20779 7986
rect 16941 7928 16946 7984
rect 17002 7928 20718 7984
rect 20774 7928 20779 7984
rect 16941 7926 20779 7928
rect 16941 7923 17007 7926
rect 20713 7923 20779 7926
rect 21449 7986 21515 7989
rect 22200 7986 23000 8016
rect 21449 7984 23000 7986
rect 21449 7928 21454 7984
rect 21510 7928 23000 7984
rect 21449 7926 23000 7928
rect 21449 7923 21515 7926
rect 22200 7896 23000 7926
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 22200 7578 23000 7608
rect 22142 7488 23000 7578
rect 21357 7442 21423 7445
rect 22142 7442 22202 7488
rect 21357 7440 22202 7442
rect 21357 7384 21362 7440
rect 21418 7384 22202 7440
rect 21357 7382 22202 7384
rect 21357 7379 21423 7382
rect 20345 7170 20411 7173
rect 22200 7170 23000 7200
rect 20345 7168 23000 7170
rect 20345 7112 20350 7168
rect 20406 7112 23000 7168
rect 20345 7110 23000 7112
rect 20345 7107 20411 7110
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 22200 7080 23000 7110
rect 19139 7039 19455 7040
rect 18086 6700 18092 6764
rect 18156 6762 18162 6764
rect 20713 6762 20779 6765
rect 18156 6760 20779 6762
rect 18156 6704 20718 6760
rect 20774 6704 20779 6760
rect 18156 6702 20779 6704
rect 18156 6700 18162 6702
rect 20713 6699 20779 6702
rect 21357 6762 21423 6765
rect 22200 6762 23000 6792
rect 21357 6760 23000 6762
rect 21357 6704 21362 6760
rect 21418 6704 23000 6760
rect 21357 6702 23000 6704
rect 21357 6699 21423 6702
rect 22200 6672 23000 6702
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 19977 6354 20043 6357
rect 22200 6354 23000 6384
rect 19977 6352 23000 6354
rect 19977 6296 19982 6352
rect 20038 6296 23000 6352
rect 19977 6294 23000 6296
rect 19977 6291 20043 6294
rect 22200 6264 23000 6294
rect 12525 6218 12591 6221
rect 20713 6218 20779 6221
rect 12525 6216 20779 6218
rect 12525 6160 12530 6216
rect 12586 6160 20718 6216
rect 20774 6160 20779 6216
rect 12525 6158 20779 6160
rect 12525 6155 12591 6158
rect 20713 6155 20779 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 22200 5946 23000 5976
rect 19566 5886 23000 5946
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 18873 5810 18939 5813
rect 19241 5810 19307 5813
rect 19566 5810 19626 5886
rect 22200 5856 23000 5886
rect 18873 5808 19626 5810
rect 18873 5752 18878 5808
rect 18934 5752 19246 5808
rect 19302 5752 19626 5808
rect 18873 5750 19626 5752
rect 18873 5747 18939 5750
rect 19241 5747 19307 5750
rect 21590 5614 22202 5674
rect 18689 5538 18755 5541
rect 20437 5538 20503 5541
rect 18689 5536 20503 5538
rect 18689 5480 18694 5536
rect 18750 5480 20442 5536
rect 20498 5480 20503 5536
rect 18689 5478 20503 5480
rect 18689 5475 18755 5478
rect 20437 5475 20503 5478
rect 20621 5538 20687 5541
rect 21590 5538 21650 5614
rect 20621 5536 21650 5538
rect 20621 5480 20626 5536
rect 20682 5480 21650 5536
rect 20621 5478 21650 5480
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 20621 5475 20687 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 11789 5130 11855 5133
rect 20345 5130 20411 5133
rect 11789 5128 20411 5130
rect 11789 5072 11794 5128
rect 11850 5072 20350 5128
rect 20406 5072 20411 5128
rect 11789 5070 20411 5072
rect 11789 5067 11855 5070
rect 20345 5067 20411 5070
rect 20621 5130 20687 5133
rect 22200 5130 23000 5160
rect 20621 5128 23000 5130
rect 20621 5072 20626 5128
rect 20682 5072 23000 5128
rect 20621 5070 23000 5072
rect 20621 5067 20687 5070
rect 22200 5040 23000 5070
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 20345 4722 20411 4725
rect 22200 4722 23000 4752
rect 20345 4720 23000 4722
rect 20345 4664 20350 4720
rect 20406 4664 23000 4720
rect 20345 4662 23000 4664
rect 20345 4659 20411 4662
rect 22200 4632 23000 4662
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 22200 4314 23000 4344
rect 22142 4224 23000 4314
rect 21357 4178 21423 4181
rect 22142 4178 22202 4224
rect 21357 4176 22202 4178
rect 21357 4120 21362 4176
rect 21418 4120 22202 4176
rect 21357 4118 22202 4120
rect 21357 4115 21423 4118
rect 20161 3906 20227 3909
rect 21265 3906 21331 3909
rect 22200 3906 23000 3936
rect 20161 3904 23000 3906
rect 20161 3848 20166 3904
rect 20222 3848 21270 3904
rect 21326 3848 23000 3904
rect 20161 3846 23000 3848
rect 20161 3843 20227 3846
rect 21265 3843 21331 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 21265 3498 21331 3501
rect 22200 3498 23000 3528
rect 21265 3496 23000 3498
rect 21265 3440 21270 3496
rect 21326 3440 23000 3496
rect 21265 3438 23000 3440
rect 21265 3435 21331 3438
rect 22200 3408 23000 3438
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 21265 3090 21331 3093
rect 22200 3090 23000 3120
rect 21265 3088 23000 3090
rect 21265 3032 21270 3088
rect 21326 3032 23000 3088
rect 21265 3030 23000 3032
rect 21265 3027 21331 3030
rect 22200 3000 23000 3030
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 20621 2682 20687 2685
rect 22200 2682 23000 2712
rect 20621 2680 23000 2682
rect 20621 2624 20626 2680
rect 20682 2624 23000 2680
rect 20621 2622 23000 2624
rect 20621 2619 20687 2622
rect 22200 2592 23000 2622
rect 20161 2410 20227 2413
rect 20161 2408 22202 2410
rect 20161 2352 20166 2408
rect 20222 2352 22202 2408
rect 20161 2350 22202 2352
rect 20161 2347 20227 2350
rect 22142 2304 22202 2350
rect 22142 2214 23000 2304
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 20253 1866 20319 1869
rect 22200 1866 23000 1896
rect 20253 1864 23000 1866
rect 20253 1808 20258 1864
rect 20314 1808 23000 1864
rect 20253 1806 23000 1808
rect 20253 1803 20319 1806
rect 22200 1776 23000 1806
rect 20529 1458 20595 1461
rect 22200 1458 23000 1488
rect 20529 1456 23000 1458
rect 20529 1400 20534 1456
rect 20590 1400 23000 1456
rect 20529 1398 23000 1400
rect 20529 1395 20595 1398
rect 22200 1368 23000 1398
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 18092 19408 18156 19412
rect 18092 19352 18106 19408
rect 18106 19352 18156 19408
rect 18092 19348 18156 19352
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 18092 6700 18156 6764
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 18091 19412 18157 19413
rect 18091 19348 18092 19412
rect 18156 19348 18157 19412
rect 18091 19347 18157 19348
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 18094 6765 18154 19347
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 18091 6764 18157 6765
rect 18091 6700 18092 6764
rect 18156 6700 18157 6764
rect 18091 6699 18157 6700
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 19872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 18584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 20792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 19688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 19320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 2024 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 7544 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 6992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 9200 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 12512 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 2208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 5336 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 4968 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 19872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 20608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8372 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_199 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1649977179
transform 1 0 20884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1649977179
transform 1 0 19872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1649977179
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_212
timestamp 1649977179
transform 1 0 20608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_216
timestamp 1649977179
transform 1 0 20976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_190
timestamp 1649977179
transform 1 0 18584 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_209
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1649977179
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1649977179
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_200
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1649977179
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1649977179
transform 1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1649977179
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1649977179
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_198
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1649977179
transform 1 0 19688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1649977179
transform 1 0 20148 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_212
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_149
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_166
timestamp 1649977179
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_178
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1649977179
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_199
timestamp 1649977179
transform 1 0 19412 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1649977179
transform 1 0 20056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_211
timestamp 1649977179
transform 1 0 20516 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_217
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_22
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_152
timestamp 1649977179
transform 1 0 15088 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_196
timestamp 1649977179
transform 1 0 19136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_201
timestamp 1649977179
transform 1 0 19596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_150
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_164
timestamp 1649977179
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_175
timestamp 1649977179
transform 1 0 17204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_217
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_123
timestamp 1649977179
transform 1 0 12420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_147
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_154
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_189
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_194
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_198
timestamp 1649977179
transform 1 0 19320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1649977179
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1649977179
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_144
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_148
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_216
timestamp 1649977179
transform 1 0 20976 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1649977179
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_183
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_208
timestamp 1649977179
transform 1 0 20240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1649977179
transform 1 0 20608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_91
timestamp 1649977179
transform 1 0 9476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_99
timestamp 1649977179
transform 1 0 10212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1649977179
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_178
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_200
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_204
timestamp 1649977179
transform 1 0 19872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_83
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_95
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_127
timestamp 1649977179
transform 1 0 12788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_139
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_151
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_156
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_185
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1649977179
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_206
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_211
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_113
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1649977179
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_164
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_168
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_191
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1649977179
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1649977179
transform 1 0 20608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_74
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_78
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_90
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_130
timestamp 1649977179
transform 1 0 13064 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1649977179
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1649977179
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1649977179
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_116
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_173
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_75
timestamp 1649977179
transform 1 0 8004 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_87
timestamp 1649977179
transform 1 0 9108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_190
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_194
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1649977179
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_63
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_114
timestamp 1649977179
transform 1 0 11592 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_162
timestamp 1649977179
transform 1 0 16008 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_211
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_216
timestamp 1649977179
transform 1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_139
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_186
timestamp 1649977179
transform 1 0 18216 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_190
timestamp 1649977179
transform 1 0 18584 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1649977179
transform 1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_214
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_95
timestamp 1649977179
transform 1 0 9844 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_116
timestamp 1649977179
transform 1 0 11776 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_167
timestamp 1649977179
transform 1 0 16468 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_185
timestamp 1649977179
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1649977179
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_70
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_79
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp 1649977179
transform 1 0 9476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_147
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_179
timestamp 1649977179
transform 1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_216
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp 1649977179
transform 1 0 7912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_123
timestamp 1649977179
transform 1 0 12420 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1649977179
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_207
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1649977179
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_129
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_133
timestamp 1649977179
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_145
timestamp 1649977179
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_177
timestamp 1649977179
transform 1 0 17388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_201
timestamp 1649977179
transform 1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1649977179
transform 1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_214
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_50
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_62
timestamp 1649977179
transform 1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_70
timestamp 1649977179
transform 1 0 7544 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_87
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_93
timestamp 1649977179
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_143
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_155
timestamp 1649977179
transform 1 0 15364 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1649977179
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 1649977179
transform 1 0 20148 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1649977179
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1649977179
transform 1 0 20976 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_60
timestamp 1649977179
transform 1 0 6624 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_70
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_90
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_102
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_127
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_153
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1649977179
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_177
timestamp 1649977179
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_188
timestamp 1649977179
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_58
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1649977179
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_95
timestamp 1649977179
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_113
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_147
timestamp 1649977179
transform 1 0 14628 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_171
timestamp 1649977179
transform 1 0 16836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_183
timestamp 1649977179
transform 1 0 17940 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1649977179
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1649977179
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_217
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1649977179
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_115
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1649977179
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_183
timestamp 1649977179
transform 1 0 17940 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_198
timestamp 1649977179
transform 1 0 19320 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_37
timestamp 1649977179
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_49
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_57
timestamp 1649977179
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_75
timestamp 1649977179
transform 1 0 8004 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1649977179
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1649977179
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_200
timestamp 1649977179
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1649977179
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_222
timestamp 1649977179
transform 1 0 21528 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1649977179
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_66
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_70
timestamp 1649977179
transform 1 0 7544 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_74
timestamp 1649977179
transform 1 0 7912 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_88
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_115
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_147
timestamp 1649977179
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1649977179
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1649977179
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_5
timestamp 1649977179
transform 1 0 1564 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1649977179
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_47
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_57
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_61
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_73
timestamp 1649977179
transform 1 0 7820 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_94
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_98
timestamp 1649977179
transform 1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1649977179
transform 1 0 11776 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_124
timestamp 1649977179
transform 1 0 12512 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1649977179
transform 1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1649977179
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_187
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1649977179
transform 1 0 19596 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_6
timestamp 1649977179
transform 1 0 1656 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_10
timestamp 1649977179
transform 1 0 2024 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_14
timestamp 1649977179
transform 1 0 2392 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_26
timestamp 1649977179
transform 1 0 3496 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_36
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_42
timestamp 1649977179
transform 1 0 4968 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_46
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_60
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_64
timestamp 1649977179
transform 1 0 6992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_68
timestamp 1649977179
transform 1 0 7360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_72
timestamp 1649977179
transform 1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1649977179
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_88
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1649977179
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1649977179
transform 1 0 12420 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_126
timestamp 1649977179
transform 1 0 12696 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1649977179
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1649977179
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_180
timestamp 1649977179
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_8
timestamp 1649977179
transform 1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_12
timestamp 1649977179
transform 1 0 2208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_17
timestamp 1649977179
transform 1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_22
timestamp 1649977179
transform 1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1649977179
transform 1 0 4048 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_38
timestamp 1649977179
transform 1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_42
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_57
timestamp 1649977179
transform 1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_68
timestamp 1649977179
transform 1 0 7360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1649977179
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1649977179
transform 1 0 9200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_111
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1649977179
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1649977179
transform 1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_150
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_155
timestamp 1649977179
transform 1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_166
timestamp 1649977179
transform 1 0 16376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1649977179
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1649977179
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_181
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_218
timestamp 1649977179
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_222
timestamp 1649977179
transform 1 0 21528 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_14
timestamp 1649977179
transform 1 0 2392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_20
timestamp 1649977179
transform 1 0 2944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_34
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_44
timestamp 1649977179
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1649977179
transform 1 0 6808 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_72
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_94
timestamp 1649977179
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_100
timestamp 1649977179
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1649977179
transform 1 0 12144 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_126
timestamp 1649977179
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_213
timestamp 1649977179
transform 1 0 20700 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1649977179
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _48_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform -1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 20516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform 1 0 20516 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 19504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 19780 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 20332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 18124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 17848 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 17664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform 1 0 19044 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _69_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 8648 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 20240 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform 1 0 20608 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 19872 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform -1 0 17204 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform -1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1649977179
transform -1 0 20976 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1649977179
transform 1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1649977179
transform -1 0 17388 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp 1649977179
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 20148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 19596 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 20148 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 20056 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 21160 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 20332 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 20516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 9384 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 2392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 2944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 4232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1649977179
transform -1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 21436 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 21436 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 19780 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18768 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11592 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13616 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9936 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15640 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11408 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11040 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11776 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11316 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12788 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14444 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14996 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17112 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16100 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14260 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16836 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19780 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21068 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21160 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14352 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16744 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19320 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21068 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19504 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_1__106 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17112 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8740 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_1__112
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_1__99
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15272 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_6.mux_l2_in_1__100
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16284 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12420 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16192 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l1_in_1__101
timestamp 1649977179
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17204 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5704 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5520 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_10.mux_l2_in_0__107
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_12.mux_l2_in_0__108
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7912 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8556 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_14.mux_l2_in_0__109
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_0__110
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19688 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6348 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_18.mux_l2_in_0__111
timestamp 1649977179
transform -1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17112 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7360 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8372 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_20.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5796 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_22.mux_l2_in_0__114
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_1__115
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17572 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_26.mux_l2_in_0__116
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7544 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16928 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_28.mux_l2_in_0__93
timestamp 1649977179
transform 1 0 7268 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6348 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_30.mux_l2_in_0__94
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_0__95
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16284 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9752 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17940 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_34.mux_l2_in_0__96
timestamp 1649977179
transform -1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13616 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_36.mux_l2_in_0__97
timestamp 1649977179
transform -1 0 12604 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_38.mux_l2_in_0__98
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4784 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4968 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_0__102
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8280 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8004 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19044 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_0__104
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_0__105
timestamp 1649977179
transform -1 0 18952 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20056 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_0__103
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17112 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output52 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 11776 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 19228 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21160 0 1 19584
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 16 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 17 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 18 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 19 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 20 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 21 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 22 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 23 nsew signal input
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 24 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 25 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 26 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 27 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 28 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 29 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 30 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 31 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 32 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 33 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 34 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 35 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 36 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 37 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 38 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 39 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 40 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 41 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 42 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 43 nsew signal tristate
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 44 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 45 nsew signal input
flabel metal2 s 7010 22200 7066 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 46 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 47 nsew signal input
flabel metal2 s 8114 22200 8170 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 48 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 49 nsew signal input
flabel metal2 s 9218 22200 9274 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 50 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 51 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 52 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 53 nsew signal input
flabel metal2 s 11426 22200 11482 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 54 nsew signal input
flabel metal2 s 1490 22200 1546 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 55 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 56 nsew signal input
flabel metal2 s 2594 22200 2650 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 57 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 58 nsew signal input
flabel metal2 s 3698 22200 3754 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 59 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 60 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 61 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 62 nsew signal input
flabel metal2 s 5906 22200 5962 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 63 nsew signal input
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 64 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 65 nsew signal tristate
flabel metal2 s 18050 22200 18106 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 66 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 67 nsew signal tristate
flabel metal2 s 19154 22200 19210 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 68 nsew signal tristate
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 69 nsew signal tristate
flabel metal2 s 20258 22200 20314 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 70 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 71 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 72 nsew signal tristate
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 73 nsew signal tristate
flabel metal2 s 22466 22200 22522 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 74 nsew signal tristate
flabel metal2 s 12530 22200 12586 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 75 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 76 nsew signal tristate
flabel metal2 s 13634 22200 13690 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 77 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 78 nsew signal tristate
flabel metal2 s 14738 22200 14794 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 79 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 80 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 81 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 82 nsew signal tristate
flabel metal2 s 16946 22200 17002 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 83 nsew signal tristate
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 84 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_11_
port 85 nsew signal input
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 right_bottom_grid_pin_13_
port 86 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 right_bottom_grid_pin_15_
port 87 nsew signal input
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 right_bottom_grid_pin_17_
port 88 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_1_
port 89 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_3_
port 90 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_5_
port 91 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_7_
port 92 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_9_
port 93 nsew signal input
flabel metal2 s 386 22200 442 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_1_
port 94 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
