* NGSPICE file created from top_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

.subckt top_tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ bottom_width_0_height_0_subtile_0__pin_reg_out_0_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ bottom_width_0_height_0_subtile_2__pin_inpad_0_ bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0] chanx_right_in_0[10]
+ chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13] chanx_right_in_0[14]
+ chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17] chanx_right_in_0[18]
+ chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20] chanx_right_in_0[21]
+ chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24] chanx_right_in_0[25]
+ chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28] chanx_right_in_0[29]
+ chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4] chanx_right_in_0[5]
+ chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8] chanx_right_in_0[9]
+ chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11] chanx_right_out_0[12]
+ chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15] chanx_right_out_0[16]
+ chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19] chanx_right_out_0[1]
+ chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22] chanx_right_out_0[23]
+ chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26] chanx_right_out_0[27]
+ chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2] chanx_right_out_0[3]
+ chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6] chanx_right_out_0[7]
+ chanx_right_out_0[8] chanx_right_out_0[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] clk0 gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk
+ prog_reset_bottom_in reset_bottom_in right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ right_width_0_height_0_subtile_0__pin_O_10_
+ right_width_0_height_0_subtile_0__pin_O_11_ right_width_0_height_0_subtile_0__pin_O_12_
+ right_width_0_height_0_subtile_0__pin_O_13_ right_width_0_height_0_subtile_0__pin_O_14_
+ right_width_0_height_0_subtile_0__pin_O_15_ right_width_0_height_0_subtile_0__pin_O_8_
+ right_width_0_height_0_subtile_0__pin_O_9_ sc_in sc_out test_enable_bottom_in top_width_0_height_0_subtile_0__pin_O_0_
+ top_width_0_height_0_subtile_0__pin_O_1_ top_width_0_height_0_subtile_0__pin_O_2_
+ top_width_0_height_0_subtile_0__pin_O_3_ top_width_0_height_0_subtile_0__pin_O_4_
+ top_width_0_height_0_subtile_0__pin_O_5_ top_width_0_height_0_subtile_0__pin_O_6_
+ top_width_0_height_0_subtile_0__pin_O_7_ top_width_0_height_0_subtile_0__pin_cin_0_
+ top_width_0_height_0_subtile_0__pin_reg_in_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.out sky130_fd_sc_hd__buf_4
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_11.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_10.mux_l2_in_3__352 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.mux_l2_in_3__352/HI
+ net352 sky130_fd_sc_hd__conb_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
X_294_ net14 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__368 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3__368/HI
+ net368 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__313
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__313/HI
+ net313 sky130_fd_sc_hd__conb_1
XFILLER_91_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_1_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__267
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__267/HI
+ net267 sky130_fd_sc_hd__conb_1
XFILLER_85_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ sb_1__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ net38 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput231 net231 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
Xoutput220 net220 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_2.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_12.mux_l3_in_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_1_ net6 cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ sb_1__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_13.mux_l3_in_0_ sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_20.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_59_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_1__8_.mem_bottom_track_33.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_35.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_1_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_2_ net43 net12 cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_12.mux_l1_in_3_ net353 net26 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk sb_1__8_.mem_right_track_52.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_13.mux_l2_in_1_ net316 net6 sb_1__8_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_1.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_3__255 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.mux_l2_in_3__255/HI
+ net255 sky130_fd_sc_hd__conb_1
XFILLER_89_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__279
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__279/HI
+ net279 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_11.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_362_ net117 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ sb_1__8_.mux_left_track_1.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_right_track_12.mux_l3_in_0_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk sb_1__8_.mem_left_track_3.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out
+ net18 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_345_ sb_1__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net307 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
X_276_ net37 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput210 net210 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput232 net232 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_2.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__290
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__290/HI
+ net290 sky130_fd_sc_hd__conb_1
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_12.mux_l2_in_1_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_328_ sb_1__8_.mux_bottom_track_51.out VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net296 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_11.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_20.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_59_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net267 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_12.mux_l1_in_2_ net12 net86 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_44.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_13.mux_l2_in_0_ net11 sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net269 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__mux2_4
Xcby_1__8_.mux_right_ipin_1.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND
+ VPWR VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_11.ccff_head
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_361_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ sb_1__8_.mux_left_track_3.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk sb_1__8_.mem_left_track_3.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out
+ net21 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_14.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_0.mux_l2_in_3_ net351 net4 sb_1__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_344_ sb_1__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
X_275_ sb_1__8_.mux_left_track_37.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput200 net200 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__8_.mem_right_track_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_12.mux_l2_in_0_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_327_ net52 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__242 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3__242/HI
+ net242 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_2.mux_l2_in_3__354 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.mux_l2_in_3__354/HI
+ net354 sky130_fd_sc_hd__conb_1
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_13.mux_l1_in_3__342 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.mux_l1_in_3__342/HI
+ net342 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_12.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_7.mux_l2_in_3_ net350 net233 sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_0.mux_l4_in_0_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sb_1__8_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_right_track_12.mux_l1_in_1_ net68 net80 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_75_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_7 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_12.mux_l1_in_3__353 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.mux_l1_in_3__353/HI
+ net353 sky130_fd_sc_hd__conb_1
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__276
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__276/HI
+ net276 sky130_fd_sc_hd__conb_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput111 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND
+ VPWR VPWR net111 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput100 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net100 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__249 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3__249/HI
+ net249 sky130_fd_sc_hd__conb_1
XFILLER_76_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_0.mux_l3_in_1_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net114 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net298 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__mux2_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_360_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
XFILLER_26_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ sb_1__8_.mux_left_track_5.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net119 net97 VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
Xsb_1__8_.mux_bottom_track_13.mux_l1_in_0_ net224 net41 sb_1__8_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_7.mux_l4_in_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_21.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_21.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_25.mux_l2_in_0_ sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_25.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk sb_1__8_.mem_left_track_3.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_35_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_37.mux_l3_in_0_ sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out
+ net24 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_45_prog_clk cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_0.mux_l2_in_2_ net21 net92 sb_1__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_343_ sb_1__8_.mux_bottom_track_21.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_274_ net35 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 net201 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
Xoutput234 net234 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.ccff_head net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__8_.mem_right_track_0.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_7.mux_l3_in_1_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_25.mux_l1_in_1_ net322 net32 sb_1__8_.mem_bottom_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_326_ net53 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_37.mux_l2_in_1_ net329 net14 sb_1__8_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_83_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_3.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
X_309_ sb_1__8_.mux_right_track_28.out VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net288 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_7.mux_l2_in_2_ net231 net229 sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_12.mux_l1_in_0_ net102 net108 sb_1__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net285 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_8 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk cbx_1__8_.cbx_1__8_.ccff_tail net237 VGND VGND VPWR VPWR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_right_track_36.mux_l3_in_0_ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput101 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xinput112 sc_in VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_7.mux_l1_in_3_ net227 bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_1__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_0.mux_l3_in_0_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_1_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__293
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__293/HI
+ net293 sky130_fd_sc_hd__conb_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_1.mux_l3_in_0_ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_290_ sb_1__8_.mux_left_track_7.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_21.mux_l1_in_1__320 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.mux_l1_in_1__320/HI
+ net320 sky130_fd_sc_hd__conb_1
XFILLER_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_1__8_.mem_bottom_track_19.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_36.mux_l2_in_1_ net357 sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk sb_1__8_.mem_left_track_1.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.out sky130_fd_sc_hd__clkbuf_2
XFILLER_12_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_0.mux_l2_in_1_ net75 net105 sb_1__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_342_ sb_1__8_.mux_bottom_track_23.out VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__283
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__283/HI
+ net283 sky130_fd_sc_hd__conb_1
X_273_ net34 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_1.mux_l2_in_1_ net314 sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput213 net213 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
Xoutput202 net202 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail net97 VGND
+ VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_59_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_7.mux_l3_in_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_36.mux_l1_in_2_ net8 net89 sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_25.mux_l1_in_0_ net222 net62 sb_1__8_.mem_bottom_track_25.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_34_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_325_ net54 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_29.mux_l1_in_3_ net344 net231 sb_1__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_37.mux_l2_in_0_ net224 sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_27.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_27.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_45_prog_clk cby_1__8_.mem_right_ipin_10.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_1.mux_l1_in_2_ net21 net23 sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_7.mux_l2_in_3__350 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.mux_l2_in_3__350/HI
+ net350 sky130_fd_sc_hd__conb_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_308_ net9 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3_ net370 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_7.mux_l2_in_1_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_44.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__362 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3__362/HI
+ net362 sky130_fd_sc_hd__conb_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_3__265 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.mux_l2_in_3__265/HI
+ net265 sky130_fd_sc_hd__conb_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_29.mux_l3_in_0_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xinput102 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput113 test_enable_bottom_in VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_8
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_4_ sb_1__8_.mux_left_track_45.out net30
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_3_ net258 net52 cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_29_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_7.mux_l1_in_2_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net88 sb_1__8_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk sb_1__8_.mem_bottom_track_9.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3_ net243 sb_1__8_.mux_left_track_45.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_right_track_36.mux_l2_in_0_ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net280 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__mux2_2
Xsb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.out sky130_fd_sc_hd__clkbuf_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_29.mux_l2_in_1_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_4_ sb_1__8_.mux_bottom_track_41.out net92 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_45_prog_clk cby_1__8_.mem_right_ipin_13.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_0.mux_l2_in_0_ net102 sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_right_track_0.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_341_ sb_1__8_.mux_bottom_track_25.out VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_272_ net62 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__286
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__286/HI
+ net286 sky130_fd_sc_hd__conb_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_1.mux_l2_in_0_ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput214 net214 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
Xoutput203 net203 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_87_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_2.mux_l4_in_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net277 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.out sky130_fd_sc_hd__buf_4
XFILLER_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_36.mux_l1_in_1_ net71 net83 sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_324_ net24 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk cby_1__8_.ccff_tail net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_29.mux_l1_in_2_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net74 sb_1__8_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__300
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__300/HI
+ net300 sky130_fd_sc_hd__conb_1
XFILLER_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_12.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_27.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_25.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_27.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_17.mux_l2_in_1__318 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.mux_l2_in_1__318/HI
+ net318 sky130_fd_sc_hd__conb_1
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_3_ net263 sb_1__8_.mux_bottom_track_45.out cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.out sky130_fd_sc_hd__buf_4
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_1.mux_l1_in_1_ net222 net219 sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_1.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_307_ net8 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_2_ net14 cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.mux_l3_in_1_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_7.mux_l2_in_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__8_.mem_right_track_44.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__272
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__272/HI
+ net272 sky130_fd_sc_hd__conb_1
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net303 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3_ net248 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_37.mux_l1_in_0_ net33 net44 sb_1__8_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_49.mux_l2_in_0_ net335 sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_49.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput114 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput103 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net103 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_2_ net86 cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_3_ net38 net7 cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_left_track_7.mux_l1_in_1_ net70 net82 sb_1__8_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_51.mux_l2_in_0_ net337 sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_51.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_7.mux_l4_in_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_53.mux_l2_in_1__349 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.mux_l2_in_1__349/HI
+ net349 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_3_ net255 net54 cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_3__253 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.mux_l2_in_3__253/HI
+ net253 sky130_fd_sc_hd__conb_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out net5
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_2_ net30 net41 cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_29.mux_l2_in_0_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_3_ sb_1__8_.mux_bottom_track_29.out net69 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_head net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_85_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_340_ sb_1__8_.mux_bottom_track_27.out VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_271_ sb_1__8_.mux_left_track_45.out VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_7.mux_l3_in_1_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3_ net363 net58 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput215 net215 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
Xoutput226 net226 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
Xoutput204 net204 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_36.mux_l1_in_0_ net105 net111 sb_1__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_323_ sb_1__8_.mux_right_track_0.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_13.mux_l4_in_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_29.mux_l1_in_1_ net66 net78 sb_1__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__284
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__284/HI
+ net284 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_12.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_0.mux_l1_in_0_ net111 net108 sb_1__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_2_ net90 sb_1__8_.mux_bottom_track_27.out cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_70_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_4_ net35 net4 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_right_track_0.mux_l2_in_3__351 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.mux_l2_in_3__351/HI
+ net351 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_1.mux_l1_in_0_ net224 net51 sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_9.mux_l2_in_1__339 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.mux_l2_in_1__339/HI
+ net339 sky130_fd_sc_hd__conb_1
X_306_ net7 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.mux_l3_in_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_36.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_13.mux_l3_in_1_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_53.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput115 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net115
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput104 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_1_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_left_track_7.mux_l1_in_0_ net59 net46 sb_1__8_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk sb_1__8_.mem_bottom_track_7.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk
+ sb_1__8_.mem_bottom_track_13.mem_out\[1\] net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_2_ net74 sb_1__8_.mux_bottom_track_39.out cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_49.mux_l1_in_0_ net222 net49 sb_1__8_.mem_bottom_track_49.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_1_ net10 cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk
+ sb_1__8_.mem_bottom_track_45.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_45.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_2_ sb_1__8_.mux_bottom_track_17.out net76 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_51.mux_l1_in_0_ net223 net50 sb_1__8_.mem_bottom_track_51.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ net60 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__296
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__296/HI
+ net296 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_7.mux_l3_in_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_5_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_2_ net27 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_1.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__275
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__275/HI
+ net275 sky130_fd_sc_hd__conb_1
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput216 net216 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
Xoutput205 net205 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput227 net227 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__367 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3__367/HI
+ net367 sky130_fd_sc_hd__conb_1
XFILLER_48_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_2_ net48 net17 cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ sb_1__8_.mux_right_track_2.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_29.mux_l1_in_0_ net44 net39 sb_1__8_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_10.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_1_ net70 cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_3_ net41 net10 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_2_prog_clk sb_1__8_.mem_left_track_21.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ sb_1__8_.mux_right_track_36.out VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net313 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net118 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_13.mux_l3_in_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_1__8_.mem_left_track_53.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__305
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__305/HI
+ net305 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_7.mux_l1_in_2_ sb_1__8_.mux_bottom_track_15.out net77 cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__247 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3__247/HI
+ net247 sky130_fd_sc_hd__conb_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_44_prog_clk cby_1__8_.mem_right_ipin_4.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_13.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_1_ net64 cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ sb_1__8_.mem_bottom_track_43.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_45.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_78_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_13.mux_l1_in_2_ sb_1__8_.mux_bottom_track_27.out net70 cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput217 net217 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
Xoutput206 net206 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput228 net228 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_19.mem_out\[1\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_19.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
X_321_ sb_1__8_.mux_right_track_4.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_19.mux_l3_in_0_ sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_19.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_0_ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__268
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__268/HI
+ net268 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_21.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_304_ net5 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_7.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_19.mux_l2_in_1_ net319 net3 sb_1__8_.mem_bottom_track_19.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_20.mux_l1_in_3_ net355 net25 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_1__8_.mem_left_track_45.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xcby_1__8_.mux_right_ipin_7.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput106 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_44_prog_clk cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk
+ sb_1__8_.mem_bottom_track_11.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_13.mux_l2_in_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_2.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_20.mux_l3_in_0_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_13.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_32_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput207 net207 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput229 net229 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_3.mux_l2_in_3_ net345 net233 sb_1__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_19.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_19.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_320_ sb_1__8_.mux_right_track_6.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_20.mux_l2_in_1_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xsb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_36.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__270
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__270/HI
+ net270 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_13.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_303_ net4 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_7.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_19.mux_l2_in_0_ net7 sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_19.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_20.mux_l1_in_2_ net11 net87 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_3.mux_l4_in_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mux_right_ipin_7.mux_l2_in_3__263 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.mux_l2_in_3__263/HI
+ net263 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_13.mux_l1_in_3_ net342 net229 sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_7.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_21.mux_l2_in_0_ sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_49.mux_l2_in_0__335 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.mux_l2_in_0__335/HI
+ net335 sky130_fd_sc_hd__conb_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput107 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net294 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_3.mux_l3_in_1_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_21.mux_l1_in_1_ net320 net5 sb_1__8_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net266 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_6.mux_l2_in_3_ net361 net29 sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_13.mux_l3_in_0_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_0.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_13.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput208 net208 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
XFILLER_95_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net299 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__mux2_4
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_3.mux_l2_in_2_ net230 net227 sb_1__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_17.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_19.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_20.mux_l2_in_0_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_13.mux_l2_in_1_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out
+ net23 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk sb_1__8_.mem_right_track_36.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_13_prog_clk cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ net237 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfrtp_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
X_302_ net32 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xsb_1__8_.mux_right_track_6.mux_l4_in_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_77_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_7.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_31.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_31.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_20.mux_l1_in_1_ net69 net81 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__266
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__266/HI
+ net266 sky130_fd_sc_hd__conb_1
XFILLER_59_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_left_track_13.mux_l1_in_2_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net86 sb_1__8_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput108 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND
+ VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_6.mux_l3_in_1_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_3.ccff_tail
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_19.mux_l1_in_0_ net219 net37 sb_1__8_.mem_bottom_track_19.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__280
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__280/HI
+ net280 sky130_fd_sc_hd__conb_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_3.mux_l3_in_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xinput90 chany_bottom_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_39_prog_clk
+ sb_1__8_.mem_bottom_track_37.mem_out\[1\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_37.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_21.mux_l1_in_0_ net220 net35 sb_1__8_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_33.mux_l2_in_0_ net327 sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_33.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_6.mux_l2_in_2_ net16 net74 sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_3.mux_l2_in_1_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net90 sb_1__8_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_6.mux_l1_in_3_ net66 net78 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_70_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_13.mux_l2_in_0_ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_15.mux_l2_in_1__317 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.mux_l2_in_1__317/HI
+ net317 sky130_fd_sc_hd__conb_1
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__278
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__278/HI
+ net278 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_28.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__310
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__310/HI
+ net310 sky130_fd_sc_hd__conb_1
XFILLER_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_301_ sb_1__8_.mux_right_track_44.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_6.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk
+ sb_1__8_.mem_bottom_track_29.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_31.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_45.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_20.mux_l1_in_0_ net103 net109 sb_1__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net283 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_13.mux_l1_in_1_ net68 net80 sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_21_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput109 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND
+ VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_1__8_.mux_right_track_44.mux_l3_in_0_ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.out sky130_fd_sc_hd__clkbuf_2
XFILLER_56_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_6.mux_l3_in_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3_ net239 net60 cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_7.mux_l3_in_0_ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput91 chany_bottom_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
Xinput80 chany_bottom_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_39_prog_clk
+ sb_1__8_.mem_bottom_track_37.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_37.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net284 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.out sky130_fd_sc_hd__clkbuf_2
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_44.mux_l2_in_1_ net359 sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_right_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_6.mux_l2_in_1_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_3_ net259 net53 cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_7.mux_l2_in_1_ net338 sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_3.mux_l2_in_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3_ net244 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net281 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__mux2_4
XFILLER_77_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_44.mux_l1_in_2_ net7 net90 sb_1__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_bottom_track_33.mux_l1_in_0_ net26 net56 sb_1__8_.mem_bottom_track_33.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_6.mux_l1_in_2_ net106 net104 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_13.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_45.mux_l2_in_0_ net333 sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_45.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_7.mux_l1_in_2_ net16 net19 sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ net30 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_7.mux_l2_in_1__338 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.mux_l2_in_1__338/HI
+ net338 sky130_fd_sc_hd__conb_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_3.mux_l1_in_1_ net72 net84 sb_1__8_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net114 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_3.mux_l4_in_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk sb_1__8_.mem_left_track_45.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 ccff_head_1 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_4_ net34 net32 cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_13.mux_l1_in_0_ net56 net42 sb_1__8_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_4.mem_out\[2\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_3_ net264 net52 cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__245 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3__245/HI
+ net245 sky130_fd_sc_hd__conb_1
XFILLER_20_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_37.mux_l3_in_0_ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput190 net190 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_2_ net29 net37 cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_3.mux_l3_in_1_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput70 chany_bottom_in[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
Xinput81 chany_bottom_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput92 chany_bottom_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_4
Xsb_1__8_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_35.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_37.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_3_ net249 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_4_ sb_1__8_.mux_bottom_track_41.out net92 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk net373 net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_44.mux_l2_in_0_ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_right_track_6.mux_l2_in_0_ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_37.mux_l2_in_1_ net346 sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_2_ net85 sb_1__8_.mux_bottom_track_37.out cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_7.mux_l2_in_0_ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_8.mux_l4_in_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_45_prog_clk cby_1__8_.mem_right_ipin_10.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_3_ net256 net52 cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_90_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_49.out sky130_fd_sc_hd__buf_4
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_2_ net26 cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_44.mux_l1_in_1_ net72 net84 sb_1__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_6.mux_l1_in_1_ net102 net100 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_13.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_37.mux_l1_in_2_ net232 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__8_.mem_left_track_37.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_7.mux_l1_in_1_ net222 net219 sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_8.mux_l3_in_1_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3_ net364 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net310 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__mux2_4
XFILLER_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_3.mux_l1_in_0_ net62 net48 sb_1__8_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_4_ sb_1__8_.mux_bottom_track_41.out net92 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_5.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
X_359_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk sb_1__8_.mem_left_track_37.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 ccff_head_2 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_3_ sb_1__8_.mux_left_track_29.out net9
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_14.mux_l4_in_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_19_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_45.mux_l1_in_0_ net220 net40 sb_1__8_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_4.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_2_ net86 cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_40 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput180 net180 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xoutput191 net191 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_1_ net6 cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_3.mux_l3_in_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_45_prog_clk cby_1__8_.mem_right_ipin_13.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew235 net238 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_16
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_14.mux_l3_in_1_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xinput71 chany_bottom_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput82 chany_bottom_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 net112 net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_2_ net14 net35 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_35.mux_l2_in_0__328 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.mux_l2_in_0__328/HI
+ net328 sky130_fd_sc_hd__conb_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_3_ sb_1__8_.mux_bottom_track_29.out net69 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net302 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_37.mux_l2_in_0_ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_1_ net65 cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_44_prog_clk cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_3__250 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.mux_l2_in_3__250/HI
+ net250 sky130_fd_sc_hd__conb_1
XFILLER_68_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_2_ net86 cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net273 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_42_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_44.mux_l1_in_0_ net106 net100 sb_1__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_28.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_6.mux_l1_in_0_ net110 net108 sb_1__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__288
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__288/HI
+ net288 sky130_fd_sc_hd__conb_1
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_11.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_left_track_37.mux_l1_in_1_ net63 net65 sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_3.mux_l1_in_2_ sb_1__8_.mux_bottom_track_19.out net75 cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_7.mux_l1_in_0_ net224 net46 sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_8.mux_l3_in_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_2_ net26 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_3_ sb_1__8_.mux_bottom_track_29.out net69 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_40_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk sb_1__8_.mem_left_track_5.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_358_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
X_289_ net51 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_3__261 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.mux_l2_in_3__261/HI
+ net261 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_57_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__8_.mem_right_track_4.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_1_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_3_ sb_1__8_.mux_left_track_29.out
+ net9 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_30 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput170 net170 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_45_prog_clk cby_1__8_.mem_right_ipin_13.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_12
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_14.mux_l3_in_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xinput72 chany_bottom_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xinput83 chany_bottom_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_1_ net4 cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_2_ sb_1__8_.mux_bottom_track_17.out net76 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_15.mux_l3_in_0_ sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_15.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__365 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3__365/HI
+ net365 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__241 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3__241/HI
+ net241 sky130_fd_sc_hd__conb_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_0_ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__8_.mux_right_ipin_2.mux_l2_in_3__258 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_2.mux_l2_in_3__258/HI
+ net258 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_1_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_2_ net41 net10 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_15.mux_l2_in_1_ net317 net31 sb_1__8_.mem_bottom_track_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk sb_1__8_.mem_right_track_28.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_37.mux_l1_in_0_ net77 net38 sb_1__8_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__8_.mux_right_ipin_3.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_44_prog_clk
+ sb_1__8_.mem_bottom_track_23.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_23.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__369 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3__369/HI
+ net369 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_2_ sb_1__8_.mux_bottom_track_17.out net76 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_1_prog_clk sb_1__8_.mem_left_track_5.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_357_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_288_ sb_1__8_.mux_left_track_11.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_49_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net292 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__mux2_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__8_.mem_right_track_2.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__295
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__295/HI
+ net295 sky130_fd_sc_hd__conb_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_47.mux_l2_in_0__334 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.mux_l2_in_0__334/HI
+ net334 sky130_fd_sc_hd__conb_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_20 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_42 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput160 net160 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_13.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew237 net98 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_16
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
Xinput73 chany_bottom_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xinput84 chany_bottom_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_5.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_10.ccff_head
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_0_ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net300 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net291 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_15_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_15.mux_l2_in_0_ net9 sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_15.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk sb_1__8_.mem_right_track_20.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_14.mux_l2_in_3__256 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.mux_l2_in_3__256/HI
+ net256 sky130_fd_sc_hd__conb_1
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_3.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_23.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_21.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_23.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk sb_1__8_.mem_left_track_37.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_77_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_1__8_.mem_left_track_3.ccff_tail
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_356_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
X_287_ sb_1__8_.mux_left_track_13.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_339_ sb_1__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out
+ net19 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_2.mux_l2_in_3_ net354 net32 sb_1__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_10 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput150 net150 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput161 net161 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
XFILLER_87_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ sb_1__8_.mem_bottom_track_29.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__8_.mem_right_ipin_12.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew238 net98 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_12
XFILLER_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
Xinput63 chany_bottom_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput85 chany_bottom_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput74 chany_bottom_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__312
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__312/HI
+ net312 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_5.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_8.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_2.mux_l4_in_0_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sb_1__8_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_9.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_13.mux_l2_in_1__316 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.mux_l2_in_1__316/HI
+ net316 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk sb_1__8_.mem_left_track_37.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_2.mux_l3_in_1_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_14.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_5.mux_l2_in_1__336 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.mux_l2_in_1__336/HI
+ net336 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mux_bottom_track_51.mux_l2_in_0__337 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.mux_l2_in_0__337/HI
+ net337 sky130_fd_sc_hd__conb_1
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_355_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_286_ net48 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\] net237 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_29_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_15.mux_l1_in_0_ net225 net39 sb_1__8_.mem_bottom_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_32_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_27.mux_l2_in_0_ sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_27.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__307
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__307/HI
+ net307 sky130_fd_sc_hd__conb_1
XFILLER_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net274 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__mux2_4
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ sb_1__8_.mux_bottom_track_31.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_21.mux_l1_in_3_ net343 net230 sb_1__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_269_ net59 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out
+ net22 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_right_track_2.mux_l2_in_2_ net18 net64 sb_1__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_64_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_22 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_44 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xoutput151 net151 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__243 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_3.mux_l2_in_3__243/HI
+ net243 sky130_fd_sc_hd__conb_1
XFILLER_87_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput173 net173 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ sb_1__8_.mem_bottom_track_27.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__303
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__303/HI
+ net303 sky130_fd_sc_hd__conb_1
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_44_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput64 chany_bottom_in[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 chany_bottom_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xinput86 chany_bottom_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_27.mux_l1_in_1_ net323 net30 sb_1__8_.mem_bottom_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_3.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net289 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_41.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk
+ sb_1__8_.mem_bottom_track_41.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_41.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_21.mux_l3_in_0_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net309 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_29.mux_l2_in_0__324 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.mux_l2_in_0__324/HI
+ net324 sky130_fd_sc_hd__conb_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_81_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_21.mux_l2_in_1_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_58_prog_clk sb_1__8_.mem_left_track_29.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_94_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_2.mux_l3_in_0_ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_354_ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_285_ net47 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.out sky130_fd_sc_hd__clkbuf_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_3.mux_l3_in_0_ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_1_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_49_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__298
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__298/HI
+ net298 sky130_fd_sc_hd__conb_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_1__8_.mux_bottom_track_33.out VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_left_track_21.mux_l1_in_2_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net85 sb_1__8_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_268_ net58 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_2.mux_l2_in_1_ net76 net106 sb_1__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_37_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_23 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.out sky130_fd_sc_hd__clkbuf_2
XFILLER_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_3.mux_l2_in_1_ net325 sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput87 chany_bottom_in[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
Xinput76 chany_bottom_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput98 prog_reset_bottom_in VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
Xinput65 chany_bottom_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_0.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_88_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_27.mux_l1_in_0_ net223 net60 sb_1__8_.mem_bottom_track_27.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_39.mux_l2_in_0_ net330 sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_39.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3_ net366 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_41.mux_l2_in_0_ net331 sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_41.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_41.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk
+ net371 net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_41.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_3.mux_l1_in_2_ net18 net22 sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_left_track_45.mux_l2_in_1__347 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.mux_l2_in_1__347/HI
+ net347 sky130_fd_sc_hd__conb_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3_ net240 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_15_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_4_ sb_1__8_.mux_left_track_45.out net30
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk
+ sb_1__8_.mem_bottom_track_15.mem_out\[1\] net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_15.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_21.mux_l2_in_0_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out net5
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_3_ net260 net54 cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_51.out sky130_fd_sc_hd__clkbuf_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_29_prog_clk
+ sb_1__8_.mem_bottom_track_47.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_47.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_353_ sb_1__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_284_ net46 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_50_prog_clk cby_1__8_.mem_right_ipin_3.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_3_ net245 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ sb_1__8_.mux_bottom_track_35.out VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_left_track_21.mux_l1_in_1_ net67 net79 sb_1__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_4_ sb_1__8_.mux_bottom_track_45.out net90 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
X_267_ sb_1__8_.mux_left_track_53.out VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_2.mux_l2_in_0_ net103 sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_13 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput120 net120 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_right_track_52.mux_l3_in_0_ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xoutput197 net197 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
XFILLER_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_20_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_3.mux_l2_in_0_ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_4.mux_l4_in_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_3_ net252 net54 cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
X_319_ net21 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput66 chany_bottom_in[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xinput88 chany_bottom_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput77 chany_bottom_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xinput99 reset_bottom_in VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_8
Xsb_1__8_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.out sky130_fd_sc_hd__buf_4
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__370 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_12.mux_l2_in_3__370/HI
+ net370 sky130_fd_sc_hd__conb_1
XFILLER_87_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_2_ net14 cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_33.mux_l2_in_0__327 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_33.mux_l2_in_0__327/HI
+ net327 sky130_fd_sc_hd__conb_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.out sky130_fd_sc_hd__clkbuf_1
XFILLER_24_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__363 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_1.mux_l2_in_3__363/HI
+ net363 sky130_fd_sc_hd__conb_1
XFILLER_78_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_3_ net265 sb_1__8_.mux_bottom_track_49.out cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_52.mux_l2_in_1_ net360 net5 sb_1__8_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_3.mux_l1_in_1_ net223 net220 sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l3_in_1_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_4_ sb_1__8_.mux_bottom_track_45.out net90 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ net237 VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_36_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_39.mux_l1_in_0_ net225 net57 sb_1__8_.mem_bottom_track_39.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_3_ net38 net7 cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_6.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_10.mux_l4_in_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ sb_1__8_.mem_bottom_track_15.mem_out\[0\] net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_15.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_44.mux_l2_in_1__359 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.mux_l2_in_1__359/HI
+ net359 sky130_fd_sc_hd__conb_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_41.mux_l1_in_0_ net218 net61 sb_1__8_.mem_bottom_track_41.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_48_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net270 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_right_track_6.mux_l2_in_3__361 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_6.mux_l2_in_3__361/HI
+ net361 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_11_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_2_ net74 cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_5.mux_l2_in_3__348 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.mux_l2_in_3__348/HI
+ net348 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_9.mux_l4_in_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_30_prog_clk
+ sb_1__8_.mem_bottom_track_45.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_47.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_352_ sb_1__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_283_ sb_1__8_.mux_left_track_21.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_3_ net257 sb_1__8_.mux_bottom_track_43.out
+ cby_1__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_10.mux_l3_in_1_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk cby_1__8_.mem_right_ipin_3.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__287
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__287/HI
+ net287 sky130_fd_sc_hd__conb_1
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_2_ net28 net39 cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_10.mux_l2_in_3_ net352 net28 sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_335_ sb_1__8_.mux_bottom_track_37.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_left_track_21.mux_l1_in_0_ net55 net41 sb_1__8_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_3_ sb_1__8_.mux_bottom_track_33.out net67 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_266_ net56 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
XANTENNA_14 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_9.mux_l3_in_1_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_47 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 chanx_right_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_3_ net365 net56 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xoutput143 net143 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net311 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__mux2_4
Xoutput165 net165 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput198 net198 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_45.mux_l3_in_0_ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_2_ net74 cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
X_318_ sb_1__8_.mux_right_track_10.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput89 chany_bottom_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
Xinput67 chany_bottom_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
Xinput78 chany_bottom_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_15.mux_l4_in_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.ccff_tail VGND
+ VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_9.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_2.mux_l1_in_0_ net100 net109 sb_1__8_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_2_ net88 sb_1__8_.mux_bottom_track_31.out cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__282
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__282/HI
+ net282 sky130_fd_sc_hd__conb_1
XFILLER_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_4_ net62 net31 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_right_track_52.mux_l2_in_0_ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_10.mux_l4_in_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_3.mux_l1_in_0_ net225 net48 sb_1__8_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_45.mux_l2_in_1_ net347 net233 sb_1__8_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l3_in_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_3_ sb_1__8_.mux_bottom_track_33.out net67 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 sb_1__8_.mem_bottom_track_39.ccff_tail VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_15.mux_l3_in_1_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_81_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_58_prog_clk
+ sb_1__8_.mem_bottom_track_13.ccff_tail net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_15.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_57_prog_clk sb_1__8_.mem_left_track_29.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_10.mux_l3_in_1_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_52.mux_l1_in_1_ net91 net73 sb_1__8_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_3__254 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.mux_l2_in_3__254/HI
+ net254 sky130_fd_sc_hd__conb_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_2
XFILLER_5_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_1_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_351_ sb_1__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_282_ net43 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_2_ net91 sb_1__8_.mux_bottom_track_31.out cby_1__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.ccff_tail net97 VGND
+ VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_10.mux_l3_in_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__8_.mem_right_ipin_3.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_1_ net8 cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xsb_1__8_.mux_right_track_10.mux_l2_in_2_ net13 net85 sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net115 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ sb_1__8_.mux_bottom_track_39.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_2_ sb_1__8_.mux_bottom_track_21.out net73 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_265_ net55 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_11.mux_l3_in_0_ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_45.mux_l2_in_0__333 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_45.mux_l2_in_0__333/HI
+ net333 sky130_fd_sc_hd__conb_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_37 sb_1__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__8_.mux_right_ipin_9.mux_l3_in_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_26 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_2_ net25 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput122 net122 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_9.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__277
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__277/HI
+ net277 sky130_fd_sc_hd__conb_1
XFILLER_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_45_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net235 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_317_ sb_1__8_.mux_right_track_12.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_1_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_27.mux_l1_in_1__323 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_27.mux_l1_in_1__323/HI
+ net323 sky130_fd_sc_hd__conb_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput68 chany_bottom_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xinput79 chany_bottom_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk net1
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_2_ net46 net15 cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_10.mux_l1_in_3_ net67 net79 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_11.mux_l2_in_1_ net315 net10 sb_1__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_1_ net68 cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_3_ net39 net8 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net117 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_45.mux_l2_in_0_ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_2_ sb_1__8_.mux_bottom_track_21.out net73 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_15.mux_l3_in_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xhold2 sb_1__8_.mem_bottom_track_5.ccff_tail VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk sb_1__8_.mem_left_track_29.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_9.mux_l1_in_2_ sb_1__8_.mux_bottom_track_19.out net75 cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_10.mux_l3_in_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_95_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_52.mux_l1_in_0_ net107 net101 sb_1__8_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_88_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_45.mux_l1_in_1_ net227 net64 sb_1__8_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ sb_1__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_281_ net42 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_1_ net68 cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk cby_1__8_.mem_right_ipin_2.ccff_tail
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net306 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_10.mux_l2_in_1_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net272 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ sb_1__8_.mux_bottom_track_41.out VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_264_ net44 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_38 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput134 net134 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail net97 VGND
+ VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_0_ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_316_ net18 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_4
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput69 chany_bottom_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net293 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__mux2_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out net21
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_right_track_10.mux_l1_in_2_ net107 net105 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_37_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_11.mux_l2_in_0_ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk
+ sb_1__8_.mem_bottom_track_33.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_33.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_9.mux_l2_in_0_ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_1_ sb_1__8_.mux_bottom_track_9.out net80 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__248 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_8.mux_l2_in_3__248/HI
+ net248 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_11.mux_l1_in_1_ net12 net221 sb_1__8_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_58_prog_clk cby_1__8_.mem_right_ipin_5.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_2_prog_clk sb_1__8_.mem_left_track_21.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_9.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_45.mux_l1_in_0_ net76 net37 sb_1__8_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_11.mux_l2_in_1__315 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.mux_l2_in_1__315/HI
+ net315 sky130_fd_sc_hd__conb_1
XFILLER_67_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ net41 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_10.mux_l2_in_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ sb_1__8_.mux_bottom_track_43.out VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_4.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__309
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__309/HI
+ net309 sky130_fd_sc_hd__conb_1
XFILLER_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk sb_1__8_.mem_right_track_0.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_28 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput124 net124 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput179 net179 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_15.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_5.mux_l2_in_3_ net348 net234 sb_1__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_86_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_315_ net17 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_5.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out net24
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_10.mux_l1_in_1_ net103 net101 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__269
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__269/HI
+ net269 sky130_fd_sc_hd__conb_1
XFILLER_77_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__8_.mem_right_ipin_8.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk
+ sb_1__8_.mem_bottom_track_31.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_33.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_1_ sb_1__8_.mux_left_track_7.out
+ net21 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_10.mux_l1_in_0_ sb_1__8_.mux_bottom_track_3.out net83 cby_1__8_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_29_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_21.mux_l1_in_3__343 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_21.mux_l1_in_3__343/HI
+ net343 sky130_fd_sc_hd__conb_1
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_11.mux_l1_in_0_ net218 net42 sb_1__8_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_5.mux_l4_in_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_9.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_23.mux_l2_in_0_ sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_23.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__292
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__292/HI
+ net292 sky130_fd_sc_hd__conb_1
XFILLER_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net295 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__301
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__301/HI
+ net301 sky130_fd_sc_hd__conb_1
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mem_bottom_track_39.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk
+ sb_1__8_.mem_bottom_track_39.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_39.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xsb_1__8_.mux_left_track_3.mux_l2_in_3__345 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_3.mux_l2_in_3__345/HI
+ net345 sky130_fd_sc_hd__conb_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_3.mux_l2_in_1__325 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_3.mux_l2_in_1__325/HI
+ net325 sky130_fd_sc_hd__conb_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_left_track_5.mux_l3_in_1_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk sb_1__8_.mem_left_track_1.mem_out\[2\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_23.mux_l1_in_1_ net321 net4 sb_1__8_.mem_bottom_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_331_ sb_1__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net290 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__8_.mem_right_track_0.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_29 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput125 net125 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_5.mux_l2_in_2_ net231 net228 sb_1__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_74_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ net16 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__sdfrtp_2
Xsb_1__8_.mux_right_track_10.mux_l1_in_0_ net111 net109 sb_1__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net275 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__mux2_4
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.mux_l1_in_0_ sb_1__8_.mux_left_track_1.out
+ net24 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_6.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_8.mux_l2_in_3__264 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_8.mux_l2_in_3__264/HI
+ net264 sky130_fd_sc_hd__conb_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_13.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_bottom_track_39.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_1__8_.mem_bottom_track_37.ccff_tail net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_39.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_20.mux_l1_in_3__355 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_20.mux_l1_in_3__355/HI
+ net355 sky130_fd_sc_hd__conb_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_5.mux_l3_in_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk sb_1__8_.mem_left_track_1.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_23.mux_l1_in_0_ net221 net34 sb_1__8_.mem_bottom_track_23.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_12.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk
+ sb_1__8_.mem_bottom_track_51.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_51.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ sb_1__8_.mux_bottom_track_47.out VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_35.mux_l2_in_0_ net328 sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_35.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk sb_1__8_.mem_right_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_19 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput137 net137 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
XFILLER_55_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_3_ net368 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_5.mux_l2_in_1_ bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ net89 sb_1__8_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_313_ sb_1__8_.mux_right_track_20.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_32_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk sb_1__8_.mem_left_track_7.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_31.mux_l2_in_0__326 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.mux_l2_in_0__326/HI
+ net326 sky130_fd_sc_hd__conb_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_38_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_3_ net250 sb_1__8_.mux_bottom_track_49.out cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_4_ net34 net32 cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_6.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net304 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__mux2_4
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_41.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.out sky130_fd_sc_hd__buf_4
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_3_ net367 net44 cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk cby_1__8_.mem_right_ipin_15.mem_out\[2\]
+ net237 VGND VGND VPWR VPWR cby_1__8_.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_10.mux_l2_in_3__252 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_10.mux_l2_in_3__252/HI
+ net252 sky130_fd_sc_hd__conb_1
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__281
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__281/HI
+ net281 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_4_ sb_1__8_.mux_bottom_track_37.out net65 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_79_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_3_ net241 net58 cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_1.mux_l2_in_3__340 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.mux_l2_in_3__340/HI
+ net340 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mux_bottom_track_9.mux_l3_in_0_ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_0.mux_l4_in_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk sb_1__8_.mem_left_track_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_40_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_12.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_30_prog_clk
+ sb_1__8_.mem_bottom_track_49.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_51.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__291
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__291/HI
+ net291 sky130_fd_sc_hd__conb_1
XFILLER_6_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net308 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk net2
+ net98 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net276 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_3_ net261 net24 cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput116 net116 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput138 net138 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_9.mux_l2_in_1_ net339 sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mem_bottom_track_9.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_2_ net26 cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_0.mux_l3_in_1_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_5.mux_l2_in_0_ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_312_ net13 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
XFILLER_6_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net279 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__311
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__311/HI
+ net311 sky130_fd_sc_hd__conb_1
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3_ net246 net55 cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_7.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_35.mux_l1_in_0_ net25 net55 sb_1__8_.mem_bottom_track_35.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_39.mux_l2_in_0__330 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_39.mux_l2_in_0__330/HI
+ net330 sky130_fd_sc_hd__conb_1
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__8_.mem_bottom_track_1.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_47.mux_l2_in_0_ net334 sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_47.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_9.mux_l1_in_2_ net13 net15 sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_2_ net88 cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_3_ sb_1__8_.mux_left_track_29.out net9
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_5.mux_l1_in_1_ net71 net83 sb_1__8_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_6.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_5.mux_l4_in_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_24_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_3_ net253 net52 cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_4_ sb_1__8_.mux_left_track_45.out net30
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_2_ net3 net34 cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk cby_1__8_.mem_right_ipin_15.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_3_ sb_1__8_.mux_bottom_track_25.out net71 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_bottom_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_5.mux_l3_in_1_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_2_ net27 net35 cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__8_.mem_bottom_track_51.ccff_tail
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__8_.mux_right_ipin_11.mux_l4_in_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__274
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__274/HI
+ net274 sky130_fd_sc_hd__conb_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__366 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_0.mux_l2_in_3__366/HI
+ net366 sky130_fd_sc_hd__conb_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_2_ net63 sb_1__8_.mux_bottom_track_41.out cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_bottom_track_43.mux_l2_in_0__332 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.mux_l2_in_0__332/HI
+ net332 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_13_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput139 net139 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xsb_1__8_.mux_bottom_track_9.mux_l2_in_0_ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_9.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_0.mux_l3_in_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_311_ net12 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_52_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__8_.mem_right_track_10.mem_out\[2\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_25.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_25.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_25.mux_l1_in_1__322 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.mux_l1_in_1__322/HI
+ net322 sky130_fd_sc_hd__conb_1
XFILLER_77_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_11.mux_l3_in_1_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_2_ net14 cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk sb_1__8_.mem_left_track_7.mem_out\[0\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_1__8_.mem_bottom_track_1.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_15_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_9.mux_l1_in_1_ net223 net220 sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_42_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_1_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_2_ net47 net16 cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__8_.mux_left_track_5.mux_l1_in_0_ net60 net47 sb_1__8_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__8_.mem_right_track_4.ccff_tail
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__304
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__304/HI
+ net304 sky130_fd_sc_hd__conb_1
XFILLER_20_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_2_ net86 sb_1__8_.mux_bottom_track_35.out cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_3_ net38 net7 cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__246 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_3__246/HI
+ net246 sky130_fd_sc_hd__conb_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net286 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__mux2_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_1_ net32 cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_bottom_track_47.mux_l1_in_0_ net221 net45 sb_1__8_.mem_bottom_track_47.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk cby_1__8_.mem_right_ipin_15.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__302
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__302/HI
+ net302 sky130_fd_sc_hd__conb_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_2_ sb_1__8_.mux_bottom_track_13.out net78 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk sb_1__8_.mem_bottom_track_7.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_94_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_1_ net4 cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_5.mux_l3_in_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__271
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__271/HI
+ net271 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.out cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_2_ net43 net12 cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_11.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_1_ net92 cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput118 net118 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
XFILLER_95_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_310_ net11 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_53.mux_l3_in_0_ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.ccff_head
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__8_.mem_right_track_10.mem_out\[1\]
+ net236 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_25.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_44_prog_clk
+ sb_1__8_.mem_bottom_track_23.ccff_tail net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_25.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net297 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_11.mux_l3_in_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk sb_1__8_.mem_left_track_5.ccff_tail
+ net235 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net312 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk sb_1__8_.mem_bottom_track_1.ccff_head
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.out sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_5.mux_l1_in_2_ sb_1__8_.mux_bottom_track_23.out net72 cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_59_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_9.mux_l1_in_0_ net225 net43 sb_1__8_.mem_bottom_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_0.mux_l2_in_0_ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_53.mux_l2_in_1_ net349 net234 sb_1__8_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_15_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_1_ net66 cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_2_ sb_1__8_.mux_left_track_21.out net13
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_14.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_1_ sb_1__8_.mux_bottom_track_7.out net81 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk sb_1__8_.mem_bottom_track_7.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_11.mux_l1_in_2_ sb_1__8_.mux_bottom_track_23.out net72 cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_1_ sb_1__8_.mux_left_track_11.out net19
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_bottom_track_17.mux_l3_in_0_ sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_bottom_track_17.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_81_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_3__251 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.mux_l2_in_3__251/HI
+ net251 sky130_fd_sc_hd__conb_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_11.mux_l2_in_3_ net341 net234 sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__8_.mux_right_ipin_5.mux_l2_in_0_ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput119 net119 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__8_.mem_right_track_10.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.ccff_tail
+ net237 VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l2_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_17.mux_l2_in_1_ net318 net27 sb_1__8_.mem_bottom_track_17.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xcby_1__8_.mux_right_ipin_5.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_10.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_3__262 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.mux_l2_in_3__262/HI
+ net262 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mux_left_track_11.mux_l4_in_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sb_1__8_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_53.mux_l2_in_0_ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mux_right_ipin_11.mux_l2_in_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_1__8_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_1_ net51 net20 cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_10.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_0.mux_l1_in_0_ sb_1__8_.mux_bottom_track_1.out net84 cby_1__8_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net268 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__mux2_4
XFILLER_79_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk net372
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk
+ sb_1__8_.mem_bottom_track_11.mem_out\[1\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_11.mux_l3_in_1_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_left_track_53.mux_l1_in_1_ net228 net92 sb_1__8_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_11.mux_l1_in_1_ sb_1__8_.mux_bottom_track_11.out net79 cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_1.mux_l2_in_3_ net340 net232 sb_1__8_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_bottom_track_43.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ sb_1__8_.mem_bottom_track_43.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_43.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_8_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_1.mux_l1_in_0_ sb_1__8_.mux_left_track_5.out net22
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_36_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__8_.mux_right_ipin_3.mux_l2_in_3__259 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_3.mux_l2_in_3__259/HI
+ net259 sky130_fd_sc_hd__conb_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_11.mux_l2_in_2_ net232 net230 sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net301 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_15.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_15.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net113 VGND
+ VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__8_.mem_right_track_10.ccff_head
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ net29 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_bottom_track_17.mux_l2_in_0_ net8 sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_17.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_1.mux_l4_in_0_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sb_1__8_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__273
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__273/HI
+ net273 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_13.ccff_tail net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_3_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_11.mux_l1_in_3_ net228 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_5.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__239 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_13.mux_l2_in_3__239/HI
+ net239 sky130_fd_sc_hd__conb_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_22_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_52.mux_l2_in_1__360 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_52.mux_l2_in_1__360/HI
+ net360 sky130_fd_sc_hd__conb_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_16_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_10_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_right_track_28.mux_l1_in_3_ net356 net14 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_47_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_6.mux_l1_in_0_ sb_1__8_.mux_left_track_3.out net23
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_6.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_1.mux_l3_in_1_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_1__8_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk cby_1__8_.mem_right_ipin_2.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk
+ sb_1__8_.mem_bottom_track_11.mem_out\[0\] net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_4.mux_l2_in_3_ net358 net30 sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_11.mux_l3_in_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_53.mux_l1_in_0_ net75 net35 sb_1__8_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_1.mux_l2_in_1__314 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_1.mux_l2_in_1__314/HI
+ net314 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mux_right_ipin_11.mux_l1_in_0_ sb_1__8_.mux_bottom_track_5.out net82 cby_1__8_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_1.mux_l2_in_2_ net229 bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mem_bottom_track_43.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_1__8_.mem_bottom_track_41.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_43.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__8_.mux_right_track_28.mux_l3_in_0_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_left_track_11.mux_l2_in_1_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_72_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__285
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__285/HI
+ net285 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk
+ sb_1__8_.mem_bottom_track_17.mem_out\[1\] net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_17.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_4.mux_l4_in_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sb_1__8_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_15.mux_l2_in_3__257 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_15.mux_l2_in_3__257/HI
+ net257 sky130_fd_sc_hd__conb_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_10_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ net28 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_28.mux_l2_in_1_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk
+ sb_1__8_.mem_bottom_track_49.mem_out\[0\] net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_49.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_11.mux_l1_in_2_ bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ net87 sb_1__8_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_23_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk cby_1__8_.mem_right_ipin_5.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_4.mux_l3_in_1_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sb_1__8_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_1.ccff_tail net236 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_50_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_28.mux_l1_in_2_ net9 net88 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_17.mux_l1_in_0_ net218 net38 sb_1__8_.mem_bottom_track_17.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_1.mux_l3_in_0_ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sb_1__8_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_29.mux_l2_in_0_ net324 sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_29.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk cby_1__8_.mem_right_ipin_2.mem_out\[1\]
+ net238 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_31.mux_l2_in_0_ net326 sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_31.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk
+ sb_1__8_.mem_bottom_track_11.ccff_head net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_4.mux_l2_in_2_ net17 net63 sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_1.mux_l2_in_1_ bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ net91 sb_1__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\] net238 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__297
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__297/HI
+ net297 sky130_fd_sc_hd__conb_1
XFILLER_20_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__294
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__294/HI
+ net294 sky130_fd_sc_hd__conb_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_11.mux_l2_in_0_ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net99 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net113 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cby_1__8_.mem_right_ipin_8.mem_out\[2\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_58_prog_clk
+ sb_1__8_.mem_bottom_track_17.mem_out\[0\] net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_17.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_0_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_4.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_5.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mux_bottom_track_37.mux_l2_in_1__329 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_37.mux_l2_in_1__329/HI
+ net329 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_297_ sb_1__8_.mux_right_track_52.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_right_track_28.mux_l2_in_0_ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_30_prog_clk
+ sb_1__8_.mem_bottom_track_47.ccff_tail net98 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_49.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cbx_1__8_.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__8_.mux_left_track_11.mux_l1_in_1_ net69 net81 sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_58_prog_clk cby_1__8_.mem_right_ipin_5.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_right_track_4.mux_l3_in_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net282 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_349_ sb_1__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_left_track_29.mux_l1_in_3__344 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_29.mux_l1_in_3__344/HI
+ net344 sky130_fd_sc_hd__conb_1
XFILLER_68_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_3_ net369 net62 cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_5.mux_l3_in_0_ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_1__8_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_28.mux_l1_in_1_ net70 net82 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_25.out sky130_fd_sc_hd__clkbuf_2
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__244 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_4.mux_l2_in_3__244/HI
+ net244 sky130_fd_sc_hd__conb_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__8_.mux_left_track_37.mux_l2_in_1__346 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_37.mux_l2_in_1__346/HI
+ net346 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_11_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_2.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__289
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__289/HI
+ net289 sky130_fd_sc_hd__conb_1
Xsb_1__8_.mux_right_track_4.mux_l2_in_1_ net65 net77 sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_3_ net251 sb_1__8_.mux_bottom_track_51.out cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_5.mux_l2_in_1_ net336 net17 sb_1__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net305 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__mux2_4
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_1.mux_l2_in_0_ net73 sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.out sky130_fd_sc_hd__clkbuf_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail net235 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mem_top_ipin_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__8_.mux_bottom_track_29.mux_l1_in_0_ net29 net59 sb_1__8_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_36.mux_l2_in_1__357 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_36.mux_l2_in_1__357/HI
+ net357 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_2 chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_3_ net242 net59 cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_bottom_track_31.mux_l1_in_0_ net28 net58 sb_1__8_.mem_bottom_track_31.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_43.mux_l2_in_0_ net332 sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__8_.mem_bottom_track_43.ccff_tail VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_41.mux_l2_in_0__331 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_41.mux_l2_in_0__331/HI
+ net331 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_8.mem_out\[1\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_58_prog_clk
+ sb_1__8_.mem_bottom_track_15.ccff_tail net235 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_17.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_1.mux_l4_in_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_23.mux_l1_in_1__321 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_23.mux_l1_in_1__321/HI
+ net321 sky130_fd_sc_hd__conb_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_296_ net26 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out net5
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__mux2_1
XFILLER_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_left_track_11.mux_l1_in_0_ net58 net43 sb_1__8_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__299
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__299/HI
+ net299 sky130_fd_sc_hd__conb_1
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_5.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_3_ net262 sb_1__8_.mux_bottom_track_49.out cby_1__8_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__8_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_26_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_348_ sb_1__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_279_ sb_1__8_.mux_left_track_29.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_2_ net31 net39 cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_1.mux_l3_in_1_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_right_track_28.mux_l1_in_0_ net104 net110 sb_1__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__308
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__308/HI
+ net308 sky130_fd_sc_hd__conb_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_3_ net247 sb_1__8_.mux_left_track_53.out
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_25_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_37_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_4_ sb_1__8_.mux_bottom_track_37.out net65 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__8_.mem_right_ipin_1.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_28.mux_l1_in_3__356 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_28.mux_l1_in_3__356/HI
+ net356 sky130_fd_sc_hd__conb_1
XFILLER_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mux_right_track_4.mux_l2_in_0_ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_85_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_2_ net87 sb_1__8_.mux_bottom_track_33.out cby_1__8_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_bottom_track_5.mux_l2_in_0_ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__8_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_42_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_47.out sky130_fd_sc_hd__clkbuf_1
Xcby_1__8_.mux_right_ipin_6.mux_l4_in_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_3_ net254 sb_1__8_.mux_bottom_track_49.out
+ cby_1__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__306
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__306/HI
+ net306 sky130_fd_sc_hd__conb_1
XANTENNA_3 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_4.mux_l1_in_1_ net107 net104 sb_1__8_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__8_.mux_bottom_track_5.mux_l1_in_1_ net20 net221 sb_1__8_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_8.mem_out\[0\]
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_6.mux_l3_in_1_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_3_ net362 net59 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__8_.mux_left_track_1.mux_l1_in_0_ net34 net51 sb_1__8_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_4_ sb_1__8_.mux_bottom_track_37.out net65 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net271 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__8_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk sb_1__8_.mem_left_track_11.mem_out\[2\]
+ net238 VGND VGND VPWR VPWR sb_1__8_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_295_ net25 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l1_in_3_ net42 net11 cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_21_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_12.mux_l4_in_0_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_1__8_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_1__8_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__8_.mux_bottom_track_43.mux_l1_in_0_ net219 net36 sb_1__8_.mem_bottom_track_43.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_43.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk cby_1__8_.mem_right_ipin_4.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__8_.mux_right_ipin_6.mux_l2_in_2_ net88 cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l1_in_4_ sb_1__8_.mux_left_track_37.out
+ net5 cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_347_ sb_1__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_278_ net39 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__8_.mux_right_ipin_1.mux_l3_in_0_ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_1__8_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l2_in_1_ net8 cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_4.mux_l2_in_3__260 VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_4.mux_l2_in_3__260/HI
+ net260 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_39_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net237 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput230 net230 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__8_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND VPWR VPWR
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l4_in_0_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_12.mux_l3_in_1_ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_1__8_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_7.mux_l2_in_2_ net26 net37 cbx_1__8_.cbx_1__8_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_24_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_38_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net278 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_10_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__8_.mux_right_ipin_6.mux_l1_in_3_ sb_1__8_.mux_bottom_track_25.out net71 cby_1__8_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__8_.mux_bottom_track_19.mux_l2_in_1__319 VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_19.mux_l2_in_1__319/HI
+ net319 sky130_fd_sc_hd__conb_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_right_track_4.mux_l2_in_3__358 VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.mux_l2_in_3__358/HI
+ net358 sky130_fd_sc_hd__conb_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_1.mux_l2_in_1_ net67 cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__8_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_11.mux_l1_in_2_ sb_1__8_.mux_left_track_13.out net18
+ cbx_1__8_.cbx_1__8_.mem_top_ipin_11.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_47_prog_clk
+ sb_1__8_.mem_bottom_track_35.mem_out\[0\] net238 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_35.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_30_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_41_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net98 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l3_in_1_ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__364 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_2.mux_l2_in_3__364/HI
+ net364 sky130_fd_sc_hd__conb_1
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__8_.mux_right_ipin_12.mux_l2_in_2_ net88 cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__8_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__240 VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_14.mux_l2_in_3__240/HI
+ net240 sky130_fd_sc_hd__conb_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net287 grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__mux2_4
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__8_.mem_right_track_52.mem_out\[1\]
+ net237 VGND VGND VPWR VPWR sb_1__8_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_4 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__8_.cbx_1__8_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__8_.cbx_1__8_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_9_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net238 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__8_.mux_right_track_4.mux_l1_in_0_ net101 net110 sb_1__8_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_left_track_11.mux_l2_in_3__341 VGND VGND VPWR VPWR sb_1__8_.mux_left_track_11.mux_l2_in_3__341/HI
+ net341 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net236 VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_1.mux_l1_in_2_ sb_1__8_.mux_bottom_track_15.out net77 cby_1__8_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__8_.mux_bottom_track_5.mux_l1_in_0_ net218 net47 sb_1__8_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__8_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk cby_1__8_.mem_right_ipin_7.ccff_tail
+ net235 VGND VGND VPWR VPWR cby_1__8_.mem_right_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__8_.mux_right_ipin_6.mux_l3_in_0_ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_1__8_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.mux_l2_in_2_ net28 cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__8_.cbx_1__8_.mem_bottom_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__8_.cbx_1__8_.mux_bottom_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__8_.mux_right_ipin_12.mux_l1_in_3_ sb_1__8_.mux_bottom_track_25.out net71 cby_1__8_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__8_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
.ends

