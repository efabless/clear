magic
tech sky130A
magscale 1 2
timestamp 1656243134
<< viali >>
rect 2605 20553 2639 20587
rect 2789 20417 2823 20451
rect 1961 20349 1995 20383
rect 2237 20349 2271 20383
rect 3065 20349 3099 20383
rect 2053 20009 2087 20043
rect 2605 20009 2639 20043
rect 4445 20009 4479 20043
rect 5549 19941 5583 19975
rect 7205 19941 7239 19975
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2789 19805 2823 19839
rect 4629 19805 4663 19839
rect 5733 19805 5767 19839
rect 7389 19805 7423 19839
rect 1501 19669 1535 19703
rect 4445 19465 4479 19499
rect 8401 19465 8435 19499
rect 1685 19329 1719 19363
rect 2237 19329 2271 19363
rect 4629 19329 4663 19363
rect 8585 19329 8619 19363
rect 2053 19193 2087 19227
rect 1501 19125 1535 19159
rect 4537 18921 4571 18955
rect 1685 18717 1719 18751
rect 4721 18717 4755 18751
rect 1501 18581 1535 18615
rect 4721 18377 4755 18411
rect 1685 18241 1719 18275
rect 4905 18241 4939 18275
rect 1501 18037 1535 18071
rect 2513 17833 2547 17867
rect 3893 17833 3927 17867
rect 6929 17833 6963 17867
rect 4629 17765 4663 17799
rect 1685 17629 1719 17663
rect 2237 17629 2271 17663
rect 2697 17629 2731 17663
rect 4077 17629 4111 17663
rect 4813 17629 4847 17663
rect 7113 17629 7147 17663
rect 21097 17629 21131 17663
rect 1501 17493 1535 17527
rect 2053 17493 2087 17527
rect 20729 17493 20763 17527
rect 21281 17493 21315 17527
rect 1961 17289 1995 17323
rect 2605 17289 2639 17323
rect 3617 17289 3651 17323
rect 7297 17289 7331 17323
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2421 17153 2455 17187
rect 3801 17153 3835 17187
rect 5181 17153 5215 17187
rect 7481 17153 7515 17187
rect 4997 17017 5031 17051
rect 1501 16949 1535 16983
rect 4261 16745 4295 16779
rect 6377 16745 6411 16779
rect 9413 16609 9447 16643
rect 9597 16609 9631 16643
rect 10517 16609 10551 16643
rect 1685 16541 1719 16575
rect 4445 16541 4479 16575
rect 6561 16541 6595 16575
rect 7205 16541 7239 16575
rect 7665 16541 7699 16575
rect 9321 16473 9355 16507
rect 9965 16473 9999 16507
rect 1501 16405 1535 16439
rect 7021 16405 7055 16439
rect 7481 16405 7515 16439
rect 8953 16405 8987 16439
rect 2513 16201 2547 16235
rect 1685 16065 1719 16099
rect 1961 16065 1995 16099
rect 2697 16065 2731 16099
rect 7757 15997 7791 16031
rect 2145 15929 2179 15963
rect 1501 15861 1535 15895
rect 1961 15657 1995 15691
rect 2421 15657 2455 15691
rect 5181 15657 5215 15691
rect 7297 15657 7331 15691
rect 4353 15589 4387 15623
rect 7941 15521 7975 15555
rect 1685 15453 1719 15487
rect 2145 15453 2179 15487
rect 2605 15453 2639 15487
rect 4537 15453 4571 15487
rect 5365 15453 5399 15487
rect 7665 15453 7699 15487
rect 1501 15317 1535 15351
rect 7757 15317 7791 15351
rect 1961 15113 1995 15147
rect 2421 15113 2455 15147
rect 3341 15113 3375 15147
rect 3801 15113 3835 15147
rect 4261 15113 4295 15147
rect 4721 15113 4755 15147
rect 5273 15113 5307 15147
rect 6929 15113 6963 15147
rect 6469 15045 6503 15079
rect 1685 14977 1719 15011
rect 2145 14977 2179 15011
rect 2605 14977 2639 15011
rect 3525 14977 3559 15011
rect 3985 14977 4019 15011
rect 4629 14977 4663 15011
rect 5641 14977 5675 15011
rect 7297 14977 7331 15011
rect 7941 14977 7975 15011
rect 4813 14909 4847 14943
rect 5733 14909 5767 14943
rect 5917 14909 5951 14943
rect 7389 14909 7423 14943
rect 7573 14909 7607 14943
rect 1501 14773 1535 14807
rect 3157 14569 3191 14603
rect 9321 14569 9355 14603
rect 5181 14501 5215 14535
rect 4445 14433 4479 14467
rect 9965 14433 9999 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 2697 14365 2731 14399
rect 3341 14365 3375 14399
rect 1501 14229 1535 14263
rect 2145 14229 2179 14263
rect 2513 14229 2547 14263
rect 3801 14229 3835 14263
rect 4169 14229 4203 14263
rect 4261 14229 4295 14263
rect 8953 14229 8987 14263
rect 9689 14229 9723 14263
rect 9781 14229 9815 14263
rect 10333 14229 10367 14263
rect 11161 14229 11195 14263
rect 12449 14229 12483 14263
rect 1961 14025 1995 14059
rect 2421 14025 2455 14059
rect 4077 14025 4111 14059
rect 4905 14025 4939 14059
rect 5917 14025 5951 14059
rect 7941 14025 7975 14059
rect 8309 14025 8343 14059
rect 9413 14025 9447 14059
rect 9781 14025 9815 14059
rect 10425 14025 10459 14059
rect 10793 14025 10827 14059
rect 11529 14025 11563 14059
rect 12541 14025 12575 14059
rect 12909 14025 12943 14059
rect 6469 13957 6503 13991
rect 7665 13957 7699 13991
rect 8953 13957 8987 13991
rect 9873 13957 9907 13991
rect 1685 13889 1719 13923
rect 2145 13889 2179 13923
rect 2605 13889 2639 13923
rect 3065 13889 3099 13923
rect 3617 13889 3651 13923
rect 3709 13889 3743 13923
rect 4353 13889 4387 13923
rect 5273 13889 5307 13923
rect 8401 13889 8435 13923
rect 10885 13889 10919 13923
rect 11897 13889 11931 13923
rect 11989 13889 12023 13923
rect 3433 13821 3467 13855
rect 5365 13821 5399 13855
rect 5549 13821 5583 13855
rect 8493 13821 8527 13855
rect 10057 13821 10091 13855
rect 11069 13821 11103 13855
rect 12173 13821 12207 13855
rect 13001 13821 13035 13855
rect 13185 13821 13219 13855
rect 1501 13685 1535 13719
rect 2881 13685 2915 13719
rect 2789 13481 2823 13515
rect 3249 13481 3283 13515
rect 4169 13481 4203 13515
rect 7757 13481 7791 13515
rect 12081 13481 12115 13515
rect 7297 13413 7331 13447
rect 11437 13413 11471 13447
rect 1961 13345 1995 13379
rect 4813 13345 4847 13379
rect 5273 13345 5307 13379
rect 6285 13345 6319 13379
rect 6469 13345 6503 13379
rect 8309 13345 8343 13379
rect 10885 13345 10919 13379
rect 11713 13345 11747 13379
rect 12725 13345 12759 13379
rect 2973 13277 3007 13311
rect 3433 13277 3467 13311
rect 4537 13277 4571 13311
rect 8125 13277 8159 13311
rect 9965 13277 9999 13311
rect 10609 13277 10643 13311
rect 6193 13209 6227 13243
rect 8217 13209 8251 13243
rect 12449 13209 12483 13243
rect 1501 13141 1535 13175
rect 2053 13141 2087 13175
rect 2145 13141 2179 13175
rect 2513 13141 2547 13175
rect 4629 13141 4663 13175
rect 5825 13141 5859 13175
rect 6929 13141 6963 13175
rect 10241 13141 10275 13175
rect 10701 13141 10735 13175
rect 12541 13141 12575 13175
rect 13093 13141 13127 13175
rect 20913 13141 20947 13175
rect 1501 12937 1535 12971
rect 1961 12937 1995 12971
rect 2421 12937 2455 12971
rect 3065 12937 3099 12971
rect 5641 12937 5675 12971
rect 7389 12937 7423 12971
rect 7849 12937 7883 12971
rect 8493 12937 8527 12971
rect 12173 12937 12207 12971
rect 12541 12937 12575 12971
rect 1685 12801 1719 12835
rect 2145 12801 2179 12835
rect 2605 12801 2639 12835
rect 3249 12801 3283 12835
rect 7757 12801 7791 12835
rect 9045 12801 9079 12835
rect 10149 12801 10183 12835
rect 5733 12733 5767 12767
rect 5825 12733 5859 12767
rect 6653 12733 6687 12767
rect 7113 12733 7147 12767
rect 7941 12733 7975 12767
rect 9505 12733 9539 12767
rect 9965 12733 9999 12767
rect 10057 12733 10091 12767
rect 12633 12733 12667 12767
rect 12817 12733 12851 12767
rect 3893 12665 3927 12699
rect 10517 12665 10551 12699
rect 20453 12665 20487 12699
rect 3525 12597 3559 12631
rect 5273 12597 5307 12631
rect 20729 12597 20763 12631
rect 21189 12597 21223 12631
rect 4353 12393 4387 12427
rect 5825 12393 5859 12427
rect 6837 12393 6871 12427
rect 9321 12393 9355 12427
rect 1593 12325 1627 12359
rect 2697 12257 2731 12291
rect 4813 12257 4847 12291
rect 4997 12257 5031 12291
rect 6469 12257 6503 12291
rect 7481 12257 7515 12291
rect 8401 12257 8435 12291
rect 9873 12257 9907 12291
rect 10977 12257 11011 12291
rect 1409 12189 1443 12223
rect 2513 12189 2547 12223
rect 3341 12189 3375 12223
rect 7205 12189 7239 12223
rect 8217 12189 8251 12223
rect 9689 12189 9723 12223
rect 11805 12189 11839 12223
rect 13461 12189 13495 12223
rect 17049 12189 17083 12223
rect 20545 12189 20579 12223
rect 2605 12121 2639 12155
rect 3801 12121 3835 12155
rect 12050 12121 12084 12155
rect 16804 12121 16838 12155
rect 19901 12121 19935 12155
rect 20269 12121 20303 12155
rect 2145 12053 2179 12087
rect 3157 12053 3191 12087
rect 4721 12053 4755 12087
rect 5365 12053 5399 12087
rect 6193 12053 6227 12087
rect 6285 12053 6319 12087
rect 7297 12053 7331 12087
rect 7849 12053 7883 12087
rect 8309 12053 8343 12087
rect 9045 12053 9079 12087
rect 9781 12053 9815 12087
rect 10333 12053 10367 12087
rect 10701 12053 10735 12087
rect 10793 12053 10827 12087
rect 13185 12053 13219 12087
rect 15669 12053 15703 12087
rect 17417 12053 17451 12087
rect 21005 12053 21039 12087
rect 21373 12053 21407 12087
rect 2513 11849 2547 11883
rect 3157 11849 3191 11883
rect 4997 11849 5031 11883
rect 5457 11849 5491 11883
rect 6377 11849 6411 11883
rect 6745 11849 6779 11883
rect 6837 11849 6871 11883
rect 7757 11849 7791 11883
rect 8217 11849 8251 11883
rect 8769 11849 8803 11883
rect 9229 11849 9263 11883
rect 9781 11849 9815 11883
rect 15577 11849 15611 11883
rect 19993 11849 20027 11883
rect 4353 11781 4387 11815
rect 5365 11781 5399 11815
rect 21106 11781 21140 11815
rect 1409 11713 1443 11747
rect 3341 11713 3375 11747
rect 4445 11713 4479 11747
rect 8125 11713 8159 11747
rect 9137 11713 9171 11747
rect 10905 11713 10939 11747
rect 12337 11713 12371 11747
rect 13829 11713 13863 11747
rect 14197 11713 14231 11747
rect 14453 11713 14487 11747
rect 15945 11713 15979 11747
rect 16313 11713 16347 11747
rect 16681 11713 16715 11747
rect 16937 11713 16971 11747
rect 18593 11713 18627 11747
rect 21373 11713 21407 11747
rect 2605 11645 2639 11679
rect 2743 11645 2777 11679
rect 4537 11645 4571 11679
rect 5641 11645 5675 11679
rect 7021 11645 7055 11679
rect 8401 11645 8435 11679
rect 9413 11645 9447 11679
rect 11161 11645 11195 11679
rect 12081 11645 12115 11679
rect 18337 11645 18371 11679
rect 3985 11577 4019 11611
rect 1593 11509 1627 11543
rect 2145 11509 2179 11543
rect 3709 11509 3743 11543
rect 11621 11509 11655 11543
rect 13461 11509 13495 11543
rect 18061 11509 18095 11543
rect 19717 11509 19751 11543
rect 1409 11305 1443 11339
rect 2513 11305 2547 11339
rect 3249 11305 3283 11339
rect 4537 11305 4571 11339
rect 12081 11305 12115 11339
rect 14473 11305 14507 11339
rect 17509 11305 17543 11339
rect 19349 11305 19383 11339
rect 21097 11305 21131 11339
rect 5549 11237 5583 11271
rect 7849 11237 7883 11271
rect 12357 11237 12391 11271
rect 1961 11169 1995 11203
rect 2053 11169 2087 11203
rect 4997 11169 5031 11203
rect 5181 11169 5215 11203
rect 6193 11169 6227 11203
rect 8401 11169 8435 11203
rect 8953 11169 8987 11203
rect 13737 11169 13771 11203
rect 14105 11169 14139 11203
rect 20729 11169 20763 11203
rect 4169 11101 4203 11135
rect 5917 11101 5951 11135
rect 7481 11101 7515 11135
rect 8217 11101 8251 11135
rect 10701 11101 10735 11135
rect 10968 11101 11002 11135
rect 15586 11101 15620 11135
rect 15853 11101 15887 11135
rect 16129 11101 16163 11135
rect 17877 11101 17911 11135
rect 18245 11101 18279 11135
rect 18613 11101 18647 11135
rect 3801 11033 3835 11067
rect 13470 11033 13504 11067
rect 16396 11033 16430 11067
rect 20462 11033 20496 11067
rect 2145 10965 2179 10999
rect 2789 10965 2823 10999
rect 4905 10965 4939 10999
rect 6009 10965 6043 10999
rect 6561 10965 6595 10999
rect 8309 10965 8343 10999
rect 1961 10761 1995 10795
rect 2421 10761 2455 10795
rect 3249 10761 3283 10795
rect 3801 10761 3835 10795
rect 4261 10761 4295 10795
rect 5457 10761 5491 10795
rect 7205 10761 7239 10795
rect 18337 10761 18371 10795
rect 2329 10693 2363 10727
rect 8953 10693 8987 10727
rect 14228 10693 14262 10727
rect 1409 10625 1443 10659
rect 3893 10625 3927 10659
rect 5089 10625 5123 10659
rect 7297 10625 7331 10659
rect 7941 10625 7975 10659
rect 8861 10625 8895 10659
rect 12265 10625 12299 10659
rect 14473 10625 14507 10659
rect 15862 10625 15896 10659
rect 17794 10625 17828 10659
rect 18061 10625 18095 10659
rect 19461 10625 19495 10659
rect 19717 10625 19751 10659
rect 21106 10625 21140 10659
rect 21373 10625 21407 10659
rect 2605 10557 2639 10591
rect 3709 10557 3743 10591
rect 4905 10557 4939 10591
rect 4997 10557 5031 10591
rect 7113 10557 7147 10591
rect 8769 10557 8803 10591
rect 16129 10557 16163 10591
rect 1593 10421 1627 10455
rect 5733 10421 5767 10455
rect 6469 10421 6503 10455
rect 7665 10421 7699 10455
rect 9321 10421 9355 10455
rect 13093 10421 13127 10455
rect 14749 10421 14783 10455
rect 16681 10421 16715 10455
rect 19993 10421 20027 10455
rect 1593 10217 1627 10251
rect 2053 10217 2087 10251
rect 6193 10217 6227 10251
rect 8953 10217 8987 10251
rect 12173 10217 12207 10251
rect 17325 10217 17359 10251
rect 21005 10217 21039 10251
rect 21373 10217 21407 10251
rect 20637 10149 20671 10183
rect 3985 10081 4019 10115
rect 5089 10081 5123 10115
rect 5641 10081 5675 10115
rect 8401 10081 8435 10115
rect 9597 10081 9631 10115
rect 18705 10081 18739 10115
rect 19257 10081 19291 10115
rect 1409 10013 1443 10047
rect 1869 10013 1903 10047
rect 2329 10013 2363 10047
rect 2789 10013 2823 10047
rect 4905 10013 4939 10047
rect 9321 10013 9355 10047
rect 10793 10013 10827 10047
rect 18438 10013 18472 10047
rect 4813 9945 4847 9979
rect 5825 9945 5859 9979
rect 8309 9945 8343 9979
rect 11060 9945 11094 9979
rect 16681 9945 16715 9979
rect 19502 9945 19536 9979
rect 2513 9877 2547 9911
rect 3341 9877 3375 9911
rect 4445 9877 4479 9911
rect 5733 9877 5767 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 7573 9877 7607 9911
rect 7849 9877 7883 9911
rect 8217 9877 8251 9911
rect 9413 9877 9447 9911
rect 9965 9877 9999 9911
rect 12541 9877 12575 9911
rect 14657 9877 14691 9911
rect 16313 9877 16347 9911
rect 17049 9877 17083 9911
rect 2697 9673 2731 9707
rect 7757 9673 7791 9707
rect 9781 9673 9815 9707
rect 19349 9673 19383 9707
rect 21373 9673 21407 9707
rect 2329 9605 2363 9639
rect 5089 9605 5123 9639
rect 6745 9605 6779 9639
rect 8401 9605 8435 9639
rect 9873 9605 9907 9639
rect 12664 9605 12698 9639
rect 15577 9605 15611 9639
rect 16313 9605 16347 9639
rect 16773 9605 16807 9639
rect 20462 9605 20496 9639
rect 1409 9537 1443 9571
rect 1869 9537 1903 9571
rect 3065 9537 3099 9571
rect 3893 9537 3927 9571
rect 4997 9537 5031 9571
rect 6837 9537 6871 9571
rect 10793 9537 10827 9571
rect 12909 9537 12943 9571
rect 13185 9537 13219 9571
rect 18162 9537 18196 9571
rect 18429 9537 18463 9571
rect 18889 9537 18923 9571
rect 20729 9537 20763 9571
rect 3985 9469 4019 9503
rect 4077 9469 4111 9503
rect 5181 9469 5215 9503
rect 6929 9469 6963 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 9965 9469 9999 9503
rect 10885 9469 10919 9503
rect 11069 9469 11103 9503
rect 1593 9401 1627 9435
rect 3525 9401 3559 9435
rect 6377 9401 6411 9435
rect 7389 9401 7423 9435
rect 10425 9401 10459 9435
rect 17049 9401 17083 9435
rect 2053 9333 2087 9367
rect 4629 9333 4663 9367
rect 5641 9333 5675 9367
rect 9413 9333 9447 9367
rect 11529 9333 11563 9367
rect 15853 9333 15887 9367
rect 3249 9129 3283 9163
rect 4261 9129 4295 9163
rect 15945 9129 15979 9163
rect 17693 9129 17727 9163
rect 18245 9129 18279 9163
rect 18521 9129 18555 9163
rect 19349 9129 19383 9163
rect 19717 9129 19751 9163
rect 1593 9061 1627 9095
rect 2697 8993 2731 9027
rect 4721 8993 4755 9027
rect 4905 8993 4939 9027
rect 6929 8993 6963 9027
rect 8033 8993 8067 9027
rect 15577 8993 15611 9027
rect 17325 8993 17359 9027
rect 21097 8993 21131 9027
rect 1409 8925 1443 8959
rect 1869 8925 1903 8959
rect 3801 8925 3835 8959
rect 4629 8925 4663 8959
rect 10894 8925 10928 8959
rect 11161 8925 11195 8959
rect 12817 8925 12851 8959
rect 13093 8925 13127 8959
rect 15310 8925 15344 8959
rect 20830 8925 20864 8959
rect 5733 8857 5767 8891
rect 6469 8857 6503 8891
rect 7849 8857 7883 8891
rect 12550 8857 12584 8891
rect 17080 8857 17114 8891
rect 2053 8789 2087 8823
rect 2789 8789 2823 8823
rect 2881 8789 2915 8823
rect 3985 8789 4019 8823
rect 5273 8789 5307 8823
rect 6101 8789 6135 8823
rect 7389 8789 7423 8823
rect 7757 8789 7791 8823
rect 8401 8789 8435 8823
rect 8953 8789 8987 8823
rect 9505 8789 9539 8823
rect 9781 8789 9815 8823
rect 11437 8789 11471 8823
rect 14197 8789 14231 8823
rect 1961 8585 1995 8619
rect 2881 8585 2915 8619
rect 5273 8585 5307 8619
rect 7481 8585 7515 8619
rect 9413 8585 9447 8619
rect 9781 8585 9815 8619
rect 11161 8585 11195 8619
rect 13369 8585 13403 8619
rect 15117 8585 15151 8619
rect 15669 8585 15703 8619
rect 16221 8585 16255 8619
rect 18061 8585 18095 8619
rect 21373 8585 21407 8619
rect 3341 8517 3375 8551
rect 5365 8517 5399 8551
rect 12826 8517 12860 8551
rect 20238 8517 20272 8551
rect 1409 8449 1443 8483
rect 4261 8449 4295 8483
rect 6837 8449 6871 8483
rect 8493 8449 8527 8483
rect 13093 8449 13127 8483
rect 14482 8449 14516 8483
rect 14749 8449 14783 8483
rect 16681 8449 16715 8483
rect 16937 8449 16971 8483
rect 18337 8449 18371 8483
rect 18593 8449 18627 8483
rect 19993 8449 20027 8483
rect 2329 8381 2363 8415
rect 4353 8381 4387 8415
rect 4445 8381 4479 8415
rect 5549 8381 5583 8415
rect 7573 8381 7607 8415
rect 7757 8381 7791 8415
rect 8585 8381 8619 8415
rect 8769 8381 8803 8415
rect 9873 8381 9907 8415
rect 10057 8381 10091 8415
rect 1593 8313 1627 8347
rect 3893 8313 3927 8347
rect 5917 8313 5951 8347
rect 7113 8313 7147 8347
rect 19717 8313 19751 8347
rect 4905 8245 4939 8279
rect 8125 8245 8159 8279
rect 11713 8245 11747 8279
rect 3801 8041 3835 8075
rect 4169 8041 4203 8075
rect 6193 8041 6227 8075
rect 7205 8041 7239 8075
rect 10057 8041 10091 8075
rect 15669 8041 15703 8075
rect 17325 8041 17359 8075
rect 17601 8041 17635 8075
rect 20637 8041 20671 8075
rect 21005 8041 21039 8075
rect 21373 8041 21407 8075
rect 5917 7973 5951 8007
rect 18521 7973 18555 8007
rect 4813 7905 4847 7939
rect 5273 7905 5307 7939
rect 5457 7905 5491 7939
rect 6561 7905 6595 7939
rect 7665 7905 7699 7939
rect 7849 7905 7883 7939
rect 9505 7905 9539 7939
rect 15945 7905 15979 7939
rect 19257 7905 19291 7939
rect 1433 7837 1467 7871
rect 1869 7837 1903 7871
rect 2329 7837 2363 7871
rect 2789 7837 2823 7871
rect 3249 7837 3283 7871
rect 4537 7837 4571 7871
rect 7573 7837 7607 7871
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 12725 7837 12759 7871
rect 13277 7837 13311 7871
rect 13645 7837 13679 7871
rect 14289 7837 14323 7871
rect 18153 7837 18187 7871
rect 5549 7769 5583 7803
rect 12480 7769 12514 7803
rect 14534 7769 14568 7803
rect 16212 7769 16246 7803
rect 19524 7769 19558 7803
rect 1593 7701 1627 7735
rect 2053 7701 2087 7735
rect 2513 7701 2547 7735
rect 4629 7701 4663 7735
rect 8217 7701 8251 7735
rect 8953 7701 8987 7735
rect 10333 7701 10367 7735
rect 10701 7701 10735 7735
rect 11345 7701 11379 7735
rect 2053 7497 2087 7531
rect 2513 7497 2547 7531
rect 3985 7497 4019 7531
rect 4445 7497 4479 7531
rect 5089 7497 5123 7531
rect 7113 7497 7147 7531
rect 7481 7497 7515 7531
rect 11529 7497 11563 7531
rect 15301 7497 15335 7531
rect 15853 7497 15887 7531
rect 16129 7497 16163 7531
rect 16681 7497 16715 7531
rect 17049 7497 17083 7531
rect 17417 7497 17451 7531
rect 19073 7497 19107 7531
rect 21189 7497 21223 7531
rect 6745 7429 6779 7463
rect 7573 7429 7607 7463
rect 20729 7429 20763 7463
rect 1409 7361 1443 7395
rect 1869 7361 1903 7395
rect 2329 7361 2363 7395
rect 2789 7361 2823 7395
rect 4077 7361 4111 7395
rect 5733 7361 5767 7395
rect 8309 7361 8343 7395
rect 11069 7361 11103 7395
rect 12642 7361 12676 7395
rect 12909 7361 12943 7395
rect 13185 7361 13219 7395
rect 13553 7361 13587 7395
rect 13921 7361 13955 7395
rect 14177 7361 14211 7395
rect 18541 7361 18575 7395
rect 18797 7361 18831 7395
rect 20186 7361 20220 7395
rect 20453 7361 20487 7395
rect 3893 7293 3927 7327
rect 4813 7293 4847 7327
rect 4997 7293 5031 7327
rect 6469 7293 6503 7327
rect 7757 7293 7791 7327
rect 8585 7293 8619 7327
rect 9413 7293 9447 7327
rect 9965 7293 9999 7327
rect 2973 7225 3007 7259
rect 1593 7157 1627 7191
rect 3341 7157 3375 7191
rect 5457 7157 5491 7191
rect 8125 7157 8159 7191
rect 8953 7157 8987 7191
rect 10241 7157 10275 7191
rect 10609 7157 10643 7191
rect 5181 6953 5215 6987
rect 8953 6953 8987 6987
rect 16405 6953 16439 6987
rect 18429 6953 18463 6987
rect 18797 6953 18831 6987
rect 19257 6953 19291 6987
rect 19625 6953 19659 6987
rect 21373 6953 21407 6987
rect 13369 6885 13403 6919
rect 2237 6817 2271 6851
rect 3893 6817 3927 6851
rect 4077 6817 4111 6851
rect 5825 6817 5859 6851
rect 6837 6817 6871 6851
rect 9597 6817 9631 6851
rect 10333 6817 10367 6851
rect 11621 6817 11655 6851
rect 11989 6817 12023 6851
rect 16037 6817 16071 6851
rect 18153 6817 18187 6851
rect 21005 6817 21039 6851
rect 1409 6749 1443 6783
rect 6653 6749 6687 6783
rect 7489 6745 7523 6779
rect 7757 6749 7791 6783
rect 9321 6749 9355 6783
rect 2421 6681 2455 6715
rect 3065 6681 3099 6715
rect 4169 6681 4203 6715
rect 4813 6681 4847 6715
rect 5549 6681 5583 6715
rect 10701 6681 10735 6715
rect 11345 6681 11379 6715
rect 12245 6681 12279 6715
rect 13737 6681 13771 6715
rect 14381 6681 14415 6715
rect 15770 6681 15804 6715
rect 17908 6681 17942 6715
rect 20738 6681 20772 6715
rect 1593 6613 1627 6647
rect 2329 6613 2363 6647
rect 2789 6613 2823 6647
rect 4537 6613 4571 6647
rect 5641 6613 5675 6647
rect 6285 6613 6319 6647
rect 6745 6613 6779 6647
rect 7297 6613 7331 6647
rect 8309 6613 8343 6647
rect 9413 6613 9447 6647
rect 9965 6613 9999 6647
rect 14657 6613 14691 6647
rect 16773 6613 16807 6647
rect 4261 6409 4295 6443
rect 5641 6409 5675 6443
rect 6469 6409 6503 6443
rect 6745 6409 6779 6443
rect 8585 6409 8619 6443
rect 9045 6409 9079 6443
rect 11529 6409 11563 6443
rect 15485 6409 15519 6443
rect 15853 6409 15887 6443
rect 18061 6409 18095 6443
rect 18337 6409 18371 6443
rect 18705 6409 18739 6443
rect 19073 6409 19107 6443
rect 20821 6409 20855 6443
rect 8677 6341 8711 6375
rect 1409 6273 1443 6307
rect 2789 6273 2823 6307
rect 3249 6273 3283 6307
rect 3617 6273 3651 6307
rect 4077 6273 4111 6307
rect 4813 6273 4847 6307
rect 7113 6273 7147 6307
rect 13010 6273 13044 6307
rect 13277 6273 13311 6307
rect 14850 6273 14884 6307
rect 15117 6273 15151 6307
rect 16681 6273 16715 6307
rect 16948 6273 16982 6307
rect 19441 6273 19475 6307
rect 19697 6273 19731 6307
rect 21373 6273 21407 6307
rect 2145 6205 2179 6239
rect 5733 6205 5767 6239
rect 5825 6205 5859 6239
rect 7205 6205 7239 6239
rect 7389 6205 7423 6239
rect 8493 6205 8527 6239
rect 9321 6205 9355 6239
rect 1593 6137 1627 6171
rect 4997 6137 5031 6171
rect 2605 6069 2639 6103
rect 3065 6069 3099 6103
rect 3801 6069 3835 6103
rect 5273 6069 5307 6103
rect 8033 6069 8067 6103
rect 9781 6069 9815 6103
rect 10149 6069 10183 6103
rect 10885 6069 10919 6103
rect 11897 6069 11931 6103
rect 13737 6069 13771 6103
rect 16313 6069 16347 6103
rect 21189 6069 21223 6103
rect 3801 5865 3835 5899
rect 5273 5865 5307 5899
rect 10793 5865 10827 5899
rect 11161 5865 11195 5899
rect 13369 5865 13403 5899
rect 15853 5865 15887 5899
rect 16221 5865 16255 5899
rect 16589 5865 16623 5899
rect 18429 5865 18463 5899
rect 19349 5865 19383 5899
rect 8953 5797 8987 5831
rect 1593 5729 1627 5763
rect 2513 5729 2547 5763
rect 4721 5729 4755 5763
rect 6101 5729 6135 5763
rect 6929 5729 6963 5763
rect 7481 5729 7515 5763
rect 9597 5729 9631 5763
rect 12817 5729 12851 5763
rect 15485 5729 15519 5763
rect 17049 5729 17083 5763
rect 20729 5729 20763 5763
rect 1777 5661 1811 5695
rect 2789 5661 2823 5695
rect 3985 5661 4019 5695
rect 7573 5661 7607 5695
rect 7665 5661 7699 5695
rect 8493 5661 8527 5695
rect 9321 5661 9355 5695
rect 17305 5661 17339 5695
rect 18705 5661 18739 5695
rect 21005 5661 21039 5695
rect 1685 5593 1719 5627
rect 6193 5593 6227 5627
rect 9413 5593 9447 5627
rect 12572 5593 12606 5627
rect 15240 5593 15274 5627
rect 20462 5593 20496 5627
rect 2145 5525 2179 5559
rect 2697 5525 2731 5559
rect 3157 5525 3191 5559
rect 4813 5525 4847 5559
rect 4905 5525 4939 5559
rect 5549 5525 5583 5559
rect 6285 5525 6319 5559
rect 6653 5525 6687 5559
rect 8033 5525 8067 5559
rect 8309 5525 8343 5559
rect 9965 5525 9999 5559
rect 11437 5525 11471 5559
rect 14105 5525 14139 5559
rect 18889 5525 18923 5559
rect 21189 5525 21223 5559
rect 1593 5321 1627 5355
rect 2605 5321 2639 5355
rect 2973 5321 3007 5355
rect 3249 5321 3283 5355
rect 3709 5321 3743 5355
rect 4721 5321 4755 5355
rect 5181 5321 5215 5355
rect 6745 5321 6779 5355
rect 9137 5321 9171 5355
rect 13277 5321 13311 5355
rect 13553 5321 13587 5355
rect 16221 5321 16255 5355
rect 19441 5321 19475 5355
rect 3617 5253 3651 5287
rect 9229 5253 9263 5287
rect 10916 5253 10950 5287
rect 16948 5253 16982 5287
rect 1409 5185 1443 5219
rect 2513 5185 2547 5219
rect 4261 5185 4295 5219
rect 5089 5185 5123 5219
rect 5733 5185 5767 5219
rect 6837 5185 6871 5219
rect 7573 5185 7607 5219
rect 11161 5185 11195 5219
rect 12642 5185 12676 5219
rect 12909 5185 12943 5219
rect 15678 5185 15712 5219
rect 15945 5185 15979 5219
rect 16681 5185 16715 5219
rect 18705 5185 18739 5219
rect 19257 5185 19291 5219
rect 20830 5185 20864 5219
rect 21097 5185 21131 5219
rect 2421 5117 2455 5151
rect 3801 5117 3835 5151
rect 5365 5117 5399 5151
rect 6929 5117 6963 5151
rect 9413 5117 9447 5151
rect 8493 5049 8527 5083
rect 11529 5049 11563 5083
rect 18337 5049 18371 5083
rect 19717 5049 19751 5083
rect 1869 4981 1903 5015
rect 4445 4981 4479 5015
rect 5917 4981 5951 5015
rect 6377 4981 6411 5015
rect 7389 4981 7423 5015
rect 8125 4981 8159 5015
rect 8769 4981 8803 5015
rect 9781 4981 9815 5015
rect 13921 4981 13955 5015
rect 14565 4981 14599 5015
rect 18061 4981 18095 5015
rect 18889 4981 18923 5015
rect 4537 4777 4571 4811
rect 12633 4777 12667 4811
rect 13001 4777 13035 4811
rect 13369 4777 13403 4811
rect 13645 4777 13679 4811
rect 19257 4777 19291 4811
rect 14749 4709 14783 4743
rect 17509 4709 17543 4743
rect 1961 4641 1995 4675
rect 2237 4641 2271 4675
rect 2697 4641 2731 4675
rect 5641 4641 5675 4675
rect 5733 4641 5767 4675
rect 7297 4641 7331 4675
rect 9597 4641 9631 4675
rect 9781 4641 9815 4675
rect 11253 4641 11287 4675
rect 20637 4641 20671 4675
rect 2881 4573 2915 4607
rect 4077 4573 4111 4607
rect 4721 4573 4755 4607
rect 5181 4573 5215 4607
rect 7665 4573 7699 4607
rect 8309 4573 8343 4607
rect 10885 4573 10919 4607
rect 14473 4573 14507 4607
rect 16129 4573 16163 4607
rect 16405 4573 16439 4607
rect 18889 4573 18923 4607
rect 20913 4573 20947 4607
rect 2789 4505 2823 4539
rect 7113 4505 7147 4539
rect 11498 4505 11532 4539
rect 15862 4505 15896 4539
rect 18622 4505 18656 4539
rect 20370 4505 20404 4539
rect 3249 4437 3283 4471
rect 4261 4437 4295 4471
rect 4997 4437 5031 4471
rect 5825 4437 5859 4471
rect 6193 4437 6227 4471
rect 6653 4437 6687 4471
rect 7021 4437 7055 4471
rect 7849 4437 7883 4471
rect 8493 4437 8527 4471
rect 9137 4437 9171 4471
rect 9505 4437 9539 4471
rect 10149 4437 10183 4471
rect 14289 4437 14323 4471
rect 16589 4437 16623 4471
rect 17049 4437 17083 4471
rect 21097 4437 21131 4471
rect 3525 4233 3559 4267
rect 8953 4233 8987 4267
rect 11713 4233 11747 4267
rect 12357 4233 12391 4267
rect 5549 4165 5583 4199
rect 9321 4165 9355 4199
rect 1961 4097 1995 4131
rect 2237 4097 2271 4131
rect 2697 4097 2731 4131
rect 3341 4097 3375 4131
rect 3801 4097 3835 4131
rect 4261 4097 4295 4131
rect 4721 4097 4755 4131
rect 6469 4097 6503 4131
rect 7389 4097 7423 4131
rect 8033 4097 8067 4131
rect 8677 4097 8711 4131
rect 10149 4097 10183 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 13746 4097 13780 4131
rect 14013 4097 14047 4131
rect 15413 4097 15447 4131
rect 15669 4097 15703 4131
rect 15945 4097 15979 4131
rect 16681 4097 16715 4131
rect 16948 4097 16982 4131
rect 19450 4097 19484 4131
rect 19717 4097 19751 4131
rect 21117 4097 21151 4131
rect 21373 4097 21407 4131
rect 5641 4029 5675 4063
rect 5825 4029 5859 4063
rect 6929 4029 6963 4063
rect 9413 4029 9447 4063
rect 9505 4029 9539 4063
rect 3985 3961 4019 3995
rect 4445 3961 4479 3995
rect 4905 3961 4939 3995
rect 5181 3961 5215 3995
rect 7573 3961 7607 3995
rect 9965 3961 9999 3995
rect 10701 3961 10735 3995
rect 12633 3961 12667 3995
rect 18337 3961 18371 3995
rect 2881 3893 2915 3927
rect 6653 3893 6687 3927
rect 8217 3893 8251 3927
rect 8493 3893 8527 3927
rect 10977 3893 11011 3927
rect 14289 3893 14323 3927
rect 16129 3893 16163 3927
rect 18061 3893 18095 3927
rect 19993 3893 20027 3927
rect 4629 3689 4663 3723
rect 5549 3689 5583 3723
rect 5825 3689 5859 3723
rect 8401 3689 8435 3723
rect 16957 3689 16991 3723
rect 5089 3621 5123 3655
rect 9321 3621 9355 3655
rect 9597 3621 9631 3655
rect 11253 3621 11287 3655
rect 14105 3621 14139 3655
rect 16589 3621 16623 3655
rect 19257 3621 19291 3655
rect 1961 3553 1995 3587
rect 3341 3553 3375 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 7665 3553 7699 3587
rect 10977 3553 11011 3587
rect 15485 3553 15519 3587
rect 18337 3553 18371 3587
rect 2237 3485 2271 3519
rect 3065 3485 3099 3519
rect 3985 3485 4019 3519
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 5365 3485 5399 3519
rect 7481 3485 7515 3519
rect 7573 3485 7607 3519
rect 8585 3485 8619 3519
rect 9137 3485 9171 3519
rect 10710 3485 10744 3519
rect 12633 3485 12667 3519
rect 12909 3485 12943 3519
rect 13553 3485 13587 3519
rect 15218 3485 15252 3519
rect 15853 3485 15887 3519
rect 16405 3485 16439 3519
rect 18613 3485 18647 3519
rect 20637 3485 20671 3519
rect 20913 3485 20947 3519
rect 12366 3417 12400 3451
rect 18092 3417 18126 3451
rect 20370 3417 20404 3451
rect 4169 3349 4203 3383
rect 6193 3349 6227 3383
rect 7113 3349 7147 3383
rect 13093 3349 13127 3383
rect 13737 3349 13771 3383
rect 16037 3349 16071 3383
rect 18797 3349 18831 3383
rect 21097 3349 21131 3383
rect 5089 3145 5123 3179
rect 5549 3145 5583 3179
rect 7021 3145 7055 3179
rect 7389 3145 7423 3179
rect 8125 3145 8159 3179
rect 8585 3145 8619 3179
rect 9045 3145 9079 3179
rect 9505 3145 9539 3179
rect 13369 3145 13403 3179
rect 15025 3145 15059 3179
rect 16681 3145 16715 3179
rect 17049 3145 17083 3179
rect 1961 3009 1995 3043
rect 3617 3009 3651 3043
rect 3893 3009 3927 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 5825 3009 5859 3043
rect 6929 3009 6963 3043
rect 7941 3009 7975 3043
rect 8401 3009 8435 3043
rect 8861 2993 8895 3027
rect 9321 3009 9355 3043
rect 10894 3009 10928 3043
rect 11161 3009 11195 3043
rect 11529 3009 11563 3043
rect 11785 3009 11819 3043
rect 13185 3009 13219 3043
rect 13737 3009 13771 3043
rect 14289 3009 14323 3043
rect 14841 3009 14875 3043
rect 15393 3009 15427 3043
rect 15945 3009 15979 3043
rect 17693 3009 17727 3043
rect 18521 3009 18555 3043
rect 18777 3009 18811 3043
rect 20177 3009 20211 3043
rect 2237 2941 2271 2975
rect 3065 2941 3099 2975
rect 3341 2941 3375 2975
rect 6745 2941 6779 2975
rect 17141 2941 17175 2975
rect 17325 2941 17359 2975
rect 20545 2941 20579 2975
rect 6009 2873 6043 2907
rect 12909 2873 12943 2907
rect 9781 2805 9815 2839
rect 13921 2805 13955 2839
rect 14473 2805 14507 2839
rect 15577 2805 15611 2839
rect 16129 2805 16163 2839
rect 17877 2805 17911 2839
rect 19901 2805 19935 2839
rect 8125 2601 8159 2635
rect 9045 2601 9079 2635
rect 21281 2601 21315 2635
rect 6009 2533 6043 2567
rect 8585 2533 8619 2567
rect 11529 2533 11563 2567
rect 14289 2533 14323 2567
rect 15393 2533 15427 2567
rect 17417 2533 17451 2567
rect 1961 2465 1995 2499
rect 2237 2465 2271 2499
rect 3341 2465 3375 2499
rect 9505 2465 9539 2499
rect 12909 2465 12943 2499
rect 18061 2465 18095 2499
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 4629 2397 4663 2431
rect 4905 2397 4939 2431
rect 5365 2397 5399 2431
rect 5825 2397 5859 2431
rect 6561 2397 6595 2431
rect 7021 2397 7055 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 8401 2397 8435 2431
rect 9689 2397 9723 2431
rect 10517 2397 10551 2431
rect 11161 2397 11195 2431
rect 12653 2397 12687 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 14657 2397 14691 2431
rect 15209 2397 15243 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 18337 2397 18371 2431
rect 19441 2397 19475 2431
rect 21097 2397 21131 2431
rect 19686 2329 19720 2363
rect 5089 2261 5123 2295
rect 5549 2261 5583 2295
rect 6745 2261 6779 2295
rect 7205 2261 7239 2295
rect 7665 2261 7699 2295
rect 9597 2261 9631 2295
rect 10057 2261 10091 2295
rect 10701 2261 10735 2295
rect 10977 2261 11011 2295
rect 13369 2261 13403 2295
rect 14841 2261 14875 2295
rect 15945 2261 15979 2295
rect 16865 2261 16899 2295
rect 20821 2261 20855 2295
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2774 20584 2780 20596
rect 2639 20556 2780 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 4430 20448 4436 20460
rect 2823 20420 4436 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 4430 20408 4436 20420
rect 4488 20408 4494 20460
rect 1854 20340 1860 20392
rect 1912 20380 1918 20392
rect 1949 20383 2007 20389
rect 1949 20380 1961 20383
rect 1912 20352 1961 20380
rect 1912 20340 1918 20352
rect 1949 20349 1961 20352
rect 1995 20349 2007 20383
rect 1949 20343 2007 20349
rect 2225 20383 2283 20389
rect 2225 20349 2237 20383
rect 2271 20380 2283 20383
rect 2958 20380 2964 20392
rect 2271 20352 2964 20380
rect 2271 20349 2283 20352
rect 2225 20343 2283 20349
rect 2958 20340 2964 20352
rect 3016 20380 3022 20392
rect 3053 20383 3111 20389
rect 3053 20380 3065 20383
rect 3016 20352 3065 20380
rect 3016 20340 3022 20352
rect 3053 20349 3065 20352
rect 3099 20349 3111 20383
rect 3053 20343 3111 20349
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 2866 20040 2872 20052
rect 2639 20012 2872 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 4430 20040 4436 20052
rect 4391 20012 4436 20040
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 5537 19975 5595 19981
rect 5537 19972 5549 19975
rect 2792 19944 5549 19972
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2792 19845 2820 19944
rect 5537 19941 5549 19944
rect 5583 19941 5595 19975
rect 5537 19935 5595 19941
rect 7193 19975 7251 19981
rect 7193 19941 7205 19975
rect 7239 19941 7251 19975
rect 7193 19935 7251 19941
rect 7208 19904 7236 19935
rect 4632 19876 7236 19904
rect 4632 19845 4660 19876
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19805 2835 19839
rect 2777 19799 2835 19805
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 5718 19836 5724 19848
rect 5679 19808 5724 19836
rect 4617 19799 4675 19805
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19836 7435 19839
rect 10410 19836 10416 19848
rect 7423 19808 10416 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 2280 19468 4445 19496
rect 2280 19456 2286 19468
rect 4433 19465 4445 19468
rect 4479 19465 4491 19499
rect 4433 19459 4491 19465
rect 5718 19456 5724 19508
rect 5776 19496 5782 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 5776 19468 8401 19496
rect 5776 19456 5782 19468
rect 8389 19465 8401 19468
rect 8435 19465 8447 19499
rect 8389 19459 8447 19465
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 1946 19360 1952 19372
rect 1719 19332 1952 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 1946 19320 1952 19332
rect 2004 19320 2010 19372
rect 2222 19360 2228 19372
rect 2183 19332 2228 19360
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 4617 19363 4675 19369
rect 4617 19329 4629 19363
rect 4663 19360 4675 19363
rect 7282 19360 7288 19372
rect 4663 19332 7288 19360
rect 4663 19329 4675 19332
rect 4617 19323 4675 19329
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 8570 19360 8576 19372
rect 8531 19332 8576 19360
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 2038 19224 2044 19236
rect 1999 19196 2044 19224
rect 2038 19184 2044 19196
rect 2096 19184 2102 19236
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 1728 18924 4537 18952
rect 1728 18912 1734 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 4525 18915 4583 18921
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 3878 18748 3884 18760
rect 1719 18720 3884 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 3878 18708 3884 18720
rect 3936 18708 3942 18760
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 5902 18748 5908 18760
rect 4755 18720 5908 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 2222 18368 2228 18420
rect 2280 18408 2286 18420
rect 4709 18411 4767 18417
rect 4709 18408 4721 18411
rect 2280 18380 4721 18408
rect 2280 18368 2286 18380
rect 4709 18377 4721 18380
rect 4755 18377 4767 18411
rect 4709 18371 4767 18377
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 7466 18272 7472 18284
rect 4939 18244 7472 18272
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 1728 17836 2513 17864
rect 1728 17824 1734 17836
rect 2501 17833 2513 17836
rect 2547 17833 2559 17867
rect 3878 17864 3884 17876
rect 3839 17836 3884 17864
rect 2501 17827 2559 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 6917 17867 6975 17873
rect 6917 17864 6929 17867
rect 5960 17836 6929 17864
rect 5960 17824 5966 17836
rect 6917 17833 6929 17836
rect 6963 17833 6975 17867
rect 6917 17827 6975 17833
rect 1946 17756 1952 17808
rect 2004 17796 2010 17808
rect 4617 17799 4675 17805
rect 4617 17796 4629 17799
rect 2004 17768 4629 17796
rect 2004 17756 2010 17768
rect 4617 17765 4629 17768
rect 4663 17765 4675 17799
rect 4617 17759 4675 17765
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 1946 17660 1952 17672
rect 1719 17632 1952 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 2240 17592 2268 17623
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 2685 17663 2743 17669
rect 2685 17660 2697 17663
rect 2648 17632 2697 17660
rect 2648 17620 2654 17632
rect 2685 17629 2697 17632
rect 2731 17629 2743 17663
rect 2685 17623 2743 17629
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 6822 17660 6828 17672
rect 4847 17632 6828 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 3602 17592 3608 17604
rect 2240 17564 3608 17592
rect 3602 17552 3608 17564
rect 3660 17552 3666 17604
rect 4080 17592 4108 17623
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 9398 17660 9404 17672
rect 7147 17632 9404 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 9398 17620 9404 17632
rect 9456 17620 9462 17672
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 20732 17632 21097 17660
rect 5994 17592 6000 17604
rect 4080 17564 6000 17592
rect 5994 17552 6000 17564
rect 6052 17552 6058 17604
rect 20732 17536 20760 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2038 17524 2044 17536
rect 1999 17496 2044 17524
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 20714 17524 20720 17536
rect 20675 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21266 17524 21272 17536
rect 21227 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2590 17320 2596 17332
rect 2551 17292 2596 17320
rect 2590 17280 2596 17292
rect 2648 17280 2654 17332
rect 3602 17320 3608 17332
rect 3563 17292 3608 17320
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 7282 17320 7288 17332
rect 7243 17292 7288 17320
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17184 3847 17187
rect 5169 17187 5227 17193
rect 3835 17156 5028 17184
rect 3835 17153 3847 17156
rect 3789 17147 3847 17153
rect 2148 17048 2176 17147
rect 2424 17116 2452 17147
rect 4154 17116 4160 17128
rect 2424 17088 4160 17116
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 4246 17048 4252 17060
rect 2148 17020 4252 17048
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 5000 17057 5028 17156
rect 5169 17153 5181 17187
rect 5215 17184 5227 17187
rect 5902 17184 5908 17196
rect 5215 17156 5908 17184
rect 5215 17153 5227 17156
rect 5169 17147 5227 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 12158 17184 12164 17196
rect 7515 17156 12164 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 4985 17051 5043 17057
rect 4985 17017 4997 17051
rect 5031 17017 5043 17051
rect 4985 17011 5043 17017
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 5994 16736 6000 16788
rect 6052 16776 6058 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 6052 16748 6377 16776
rect 6052 16736 6058 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 6365 16739 6423 16745
rect 12066 16708 12072 16720
rect 9416 16680 12072 16708
rect 9416 16649 9444 16680
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16609 9459 16643
rect 9401 16603 9459 16609
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16640 9643 16643
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 9631 16612 10517 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 10505 16609 10517 16612
rect 10551 16640 10563 16643
rect 20714 16640 20720 16652
rect 10551 16612 20720 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 20714 16600 20720 16612
rect 20772 16640 20778 16652
rect 21174 16640 21180 16652
rect 20772 16612 21180 16640
rect 20772 16600 20778 16612
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2406 16572 2412 16584
rect 1719 16544 2412 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16541 4491 16575
rect 6546 16572 6552 16584
rect 6507 16544 6552 16572
rect 4433 16535 4491 16541
rect 4448 16504 4476 16535
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 7190 16572 7196 16584
rect 7151 16544 7196 16572
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 7653 16575 7711 16581
rect 7653 16541 7665 16575
rect 7699 16572 7711 16575
rect 8478 16572 8484 16584
rect 7699 16544 8484 16572
rect 7699 16541 7711 16544
rect 7653 16535 7711 16541
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 6914 16504 6920 16516
rect 4448 16476 6920 16504
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 9953 16507 10011 16513
rect 9953 16504 9965 16507
rect 9355 16476 9965 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9953 16473 9965 16476
rect 9999 16473 10011 16507
rect 9953 16467 10011 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6880 16408 7021 16436
rect 6880 16396 6886 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7466 16436 7472 16448
rect 7427 16408 7472 16436
rect 7009 16399 7067 16405
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 8570 16396 8576 16448
rect 8628 16436 8634 16448
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8628 16408 8953 16436
rect 8628 16396 8634 16408
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 1728 16204 2513 16232
rect 1728 16192 1734 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 2501 16195 2559 16201
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1946 16096 1952 16108
rect 1907 16068 1952 16096
rect 1673 16059 1731 16065
rect 1688 16028 1716 16059
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 5166 16096 5172 16108
rect 2731 16068 5172 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 2314 16028 2320 16040
rect 1688 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 7650 15988 7656 16040
rect 7708 16028 7714 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7708 16000 7757 16028
rect 7708 15988 7714 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 2130 15960 2136 15972
rect 2091 15932 2136 15960
rect 2130 15920 2136 15932
rect 2188 15920 2194 15972
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2406 15688 2412 15700
rect 2367 15660 2412 15688
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 5960 15660 7297 15688
rect 5960 15648 5966 15660
rect 7285 15657 7297 15660
rect 7331 15657 7343 15691
rect 7285 15651 7343 15657
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 2746 15592 4353 15620
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 2746 15484 2774 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 4341 15583 4399 15589
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 12250 15552 12256 15564
rect 7975 15524 12256 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 2639 15456 2774 15484
rect 4525 15487 4583 15493
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 4525 15453 4537 15487
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 5353 15487 5411 15493
rect 5353 15453 5365 15487
rect 5399 15484 5411 15487
rect 7466 15484 7472 15496
rect 5399 15456 7472 15484
rect 5399 15453 5411 15456
rect 5353 15447 5411 15453
rect 2148 15416 2176 15447
rect 3786 15416 3792 15428
rect 2148 15388 3792 15416
rect 3786 15376 3792 15388
rect 3844 15376 3850 15428
rect 4540 15416 4568 15447
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 7650 15484 7656 15496
rect 7611 15456 7656 15484
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 5994 15416 6000 15428
rect 4540 15388 6000 15416
rect 5994 15376 6000 15388
rect 6052 15376 6058 15428
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 7745 15351 7803 15357
rect 7745 15317 7757 15351
rect 7791 15348 7803 15351
rect 9306 15348 9312 15360
rect 7791 15320 9312 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1728 15116 1961 15144
rect 1728 15104 1734 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 2314 15104 2320 15156
rect 2372 15144 2378 15156
rect 2409 15147 2467 15153
rect 2409 15144 2421 15147
rect 2372 15116 2421 15144
rect 2372 15104 2378 15116
rect 2409 15113 2421 15116
rect 2455 15113 2467 15147
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 2409 15107 2467 15113
rect 2746 15116 3341 15144
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 14977 1731 15011
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 1673 14971 1731 14977
rect 1688 14940 1716 14971
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 15008 2651 15011
rect 2746 15008 2774 15116
rect 3329 15113 3341 15116
rect 3375 15113 3387 15147
rect 3786 15144 3792 15156
rect 3747 15116 3792 15144
rect 3329 15107 3387 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 4212 15116 4261 15144
rect 4212 15104 4218 15116
rect 4249 15113 4261 15116
rect 4295 15113 4307 15147
rect 4249 15107 4307 15113
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 5261 15147 5319 15153
rect 5261 15144 5273 15147
rect 4755 15116 5273 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 5261 15113 5273 15116
rect 5307 15113 5319 15147
rect 6914 15144 6920 15156
rect 6875 15116 6920 15144
rect 5261 15107 5319 15113
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 6457 15079 6515 15085
rect 6457 15076 6469 15079
rect 3988 15048 5856 15076
rect 3988 15017 4016 15048
rect 2639 14980 2774 15008
rect 3513 15011 3571 15017
rect 2639 14977 2651 14980
rect 2593 14971 2651 14977
rect 3513 14977 3525 15011
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 15008 4675 15011
rect 4890 15008 4896 15020
rect 4663 14980 4896 15008
rect 4663 14977 4675 14980
rect 4617 14971 4675 14977
rect 2406 14940 2412 14952
rect 1688 14912 2412 14940
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 3528 14872 3556 14971
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 5626 15008 5632 15020
rect 5587 14980 5632 15008
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 4798 14940 4804 14952
rect 4759 14912 4804 14940
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 5718 14940 5724 14952
rect 5679 14912 5724 14940
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 5166 14872 5172 14884
rect 3528 14844 5172 14872
rect 5166 14832 5172 14844
rect 5224 14832 5230 14884
rect 5828 14872 5856 15048
rect 5920 15048 6469 15076
rect 5920 14952 5948 15048
rect 6457 15045 6469 15048
rect 6503 15076 6515 15079
rect 15378 15076 15384 15088
rect 6503 15048 15384 15076
rect 6503 15045 6515 15048
rect 6457 15039 6515 15045
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 15008 7343 15011
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7331 14980 7941 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 7374 14940 7380 14952
rect 5960 14912 6053 14940
rect 7335 14912 7380 14940
rect 5960 14900 5966 14912
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7561 14943 7619 14949
rect 7561 14909 7573 14943
rect 7607 14909 7619 14943
rect 15562 14940 15568 14952
rect 7561 14903 7619 14909
rect 12406 14912 15568 14940
rect 7006 14872 7012 14884
rect 5828 14844 7012 14872
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 7576 14872 7604 14903
rect 12406 14872 12434 14912
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 7576 14844 12434 14872
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 2130 14560 2136 14612
rect 2188 14600 2194 14612
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 2188 14572 3157 14600
rect 2188 14560 2194 14572
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 9306 14600 9312 14612
rect 9267 14572 9312 14600
rect 3145 14563 3203 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 11698 14600 11704 14612
rect 9732 14572 11704 14600
rect 9732 14560 9738 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 13262 14600 13268 14612
rect 12406 14572 13268 14600
rect 4798 14492 4804 14544
rect 4856 14532 4862 14544
rect 5169 14535 5227 14541
rect 5169 14532 5181 14535
rect 4856 14504 5181 14532
rect 4856 14492 4862 14504
rect 5169 14501 5181 14504
rect 5215 14532 5227 14535
rect 12406 14532 12434 14572
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 5215 14504 12434 14532
rect 5215 14501 5227 14504
rect 5169 14495 5227 14501
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 9953 14467 10011 14473
rect 4479 14436 7420 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 7098 14396 7104 14408
rect 3375 14368 7104 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 2700 14328 2728 14359
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7392 14396 7420 14436
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10870 14464 10876 14476
rect 9999 14436 10876 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 10502 14396 10508 14408
rect 7392 14368 10508 14396
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 2700 14300 3832 14328
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2130 14260 2136 14272
rect 2091 14232 2136 14260
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 2501 14263 2559 14269
rect 2501 14229 2513 14263
rect 2547 14260 2559 14263
rect 2590 14260 2596 14272
rect 2547 14232 2596 14260
rect 2547 14229 2559 14232
rect 2501 14223 2559 14229
rect 2590 14220 2596 14232
rect 2648 14220 2654 14272
rect 3804 14269 3832 14300
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4028 14300 8248 14328
rect 4028 14288 4034 14300
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4157 14263 4215 14269
rect 4157 14260 4169 14263
rect 4120 14232 4169 14260
rect 4120 14220 4126 14232
rect 4157 14229 4169 14232
rect 4203 14229 4215 14263
rect 4157 14223 4215 14229
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 8220 14260 8248 14300
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 8352 14300 12480 14328
rect 8352 14288 8358 14300
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 4304 14232 4349 14260
rect 8220 14232 8953 14260
rect 4304 14220 4310 14232
rect 8941 14229 8953 14232
rect 8987 14260 8999 14263
rect 9674 14260 9680 14272
rect 8987 14232 9680 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 10318 14260 10324 14272
rect 9824 14232 9869 14260
rect 10279 14232 10324 14260
rect 9824 14220 9830 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 12452 14269 12480 14300
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10836 14232 11161 14260
rect 10836 14220 10842 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 12437 14263 12495 14269
rect 12437 14229 12449 14263
rect 12483 14260 12495 14263
rect 12894 14260 12900 14272
rect 12483 14232 12900 14260
rect 12483 14229 12495 14232
rect 12437 14223 12495 14229
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4890 14056 4896 14068
rect 4851 14028 4896 14056
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 5902 14056 5908 14068
rect 5863 14028 5908 14056
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7432 14028 7941 14056
rect 7432 14016 7438 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 8294 14056 8300 14068
rect 7929 14019 7987 14025
rect 8036 14028 8300 14056
rect 2774 13988 2780 14000
rect 1688 13960 2780 13988
rect 1688 13929 1716 13960
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 6270 13948 6276 14000
rect 6328 13988 6334 14000
rect 6457 13991 6515 13997
rect 6457 13988 6469 13991
rect 6328 13960 6469 13988
rect 6328 13948 6334 13960
rect 6457 13957 6469 13960
rect 6503 13988 6515 13991
rect 7653 13991 7711 13997
rect 7653 13988 7665 13991
rect 6503 13960 7665 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 7653 13957 7665 13960
rect 7699 13988 7711 13991
rect 8036 13988 8064 14028
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 9398 14056 9404 14068
rect 9359 14028 9404 14056
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 10318 14056 10324 14068
rect 9815 14028 10324 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 10778 14056 10784 14068
rect 10468 14028 10513 14056
rect 10739 14028 10784 14056
rect 10468 14016 10474 14028
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14025 11575 14059
rect 12529 14059 12587 14065
rect 12529 14056 12541 14059
rect 11517 14019 11575 14025
rect 11624 14028 12541 14056
rect 7699 13960 8064 13988
rect 7699 13957 7711 13960
rect 7653 13951 7711 13957
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 8941 13991 8999 13997
rect 8941 13988 8953 13991
rect 8168 13960 8953 13988
rect 8168 13948 8174 13960
rect 8941 13957 8953 13960
rect 8987 13957 8999 13991
rect 8941 13951 8999 13957
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13988 9919 13991
rect 11532 13988 11560 14019
rect 9907 13960 11560 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2133 13883 2191 13889
rect 2148 13852 2176 13883
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3384 13892 3617 13920
rect 3384 13880 3390 13892
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13920 3755 13923
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 3743 13892 4353 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 5258 13920 5264 13932
rect 5219 13892 5264 13920
rect 4341 13883 4399 13889
rect 3234 13852 3240 13864
rect 2148 13824 3240 13852
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13821 3479 13855
rect 3620 13852 3648 13883
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13920 8447 13923
rect 10873 13923 10931 13929
rect 8435 13892 10824 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 5350 13852 5356 13864
rect 3620 13824 5356 13852
rect 3421 13815 3479 13821
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 3142 13784 3148 13796
rect 1912 13756 3148 13784
rect 1912 13744 1918 13756
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 2866 13716 2872 13728
rect 2827 13688 2872 13716
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 3436 13716 3464 13815
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 5902 13852 5908 13864
rect 5583 13824 5908 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 8481 13855 8539 13861
rect 8481 13821 8493 13855
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10796 13852 10824 13892
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 11624 13920 11652 14028
rect 12529 14025 12541 14028
rect 12575 14025 12587 14059
rect 12894 14056 12900 14068
rect 12855 14028 12900 14056
rect 12529 14019 12587 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 11882 13920 11888 13932
rect 10919 13892 11652 13920
rect 11843 13892 11888 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12032 13892 12077 13920
rect 13096 13892 13308 13920
rect 12032 13880 12038 13892
rect 10962 13852 10968 13864
rect 10091 13824 10180 13852
rect 10796 13824 10968 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 8496 13784 8524 13815
rect 10152 13796 10180 13824
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 8570 13784 8576 13796
rect 8496 13756 8576 13784
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 10134 13744 10140 13796
rect 10192 13744 10198 13796
rect 4890 13716 4896 13728
rect 3436 13688 4896 13716
rect 4890 13676 4896 13688
rect 4948 13676 4954 13728
rect 11072 13716 11100 13815
rect 11146 13812 11152 13864
rect 11204 13852 11210 13864
rect 12161 13855 12219 13861
rect 11204 13824 12020 13852
rect 11204 13812 11210 13824
rect 11992 13796 12020 13824
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 11974 13744 11980 13796
rect 12032 13744 12038 13796
rect 12176 13784 12204 13815
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12400 13824 13001 13852
rect 12400 13812 12406 13824
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 13096 13784 13124 13892
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 12176 13756 13124 13784
rect 12986 13716 12992 13728
rect 11072 13688 12992 13716
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 13188 13716 13216 13815
rect 13280 13784 13308 13892
rect 13280 13756 16574 13784
rect 15654 13716 15660 13728
rect 13188 13688 15660 13716
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 16546 13716 16574 13756
rect 18966 13716 18972 13728
rect 16546 13688 18972 13716
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3234 13512 3240 13524
rect 2832 13484 2877 13512
rect 3195 13484 3240 13512
rect 2832 13472 2838 13484
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 4246 13512 4252 13524
rect 4203 13484 4252 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7248 13484 7757 13512
rect 7248 13472 7254 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 7745 13475 7803 13481
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 11790 13512 11796 13524
rect 8628 13484 11796 13512
rect 8628 13472 8634 13484
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 12066 13512 12072 13524
rect 12027 13484 12072 13512
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 7285 13447 7343 13453
rect 2746 13416 6316 13444
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 2590 13376 2596 13388
rect 1995 13348 2596 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 2746 13308 2774 13416
rect 6288 13388 6316 13416
rect 7285 13413 7297 13447
rect 7331 13444 7343 13447
rect 7834 13444 7840 13456
rect 7331 13416 7840 13444
rect 7331 13413 7343 13416
rect 7285 13407 7343 13413
rect 7834 13404 7840 13416
rect 7892 13444 7898 13456
rect 7892 13416 9996 13444
rect 7892 13404 7898 13416
rect 3142 13336 3148 13388
rect 3200 13376 3206 13388
rect 4801 13379 4859 13385
rect 3200 13348 4568 13376
rect 3200 13336 3206 13348
rect 2958 13308 2964 13320
rect 2056 13280 2774 13308
rect 2919 13280 2964 13308
rect 1489 13175 1547 13181
rect 1489 13141 1501 13175
rect 1535 13172 1547 13175
rect 1762 13172 1768 13184
rect 1535 13144 1768 13172
rect 1535 13141 1547 13144
rect 1489 13135 1547 13141
rect 1762 13132 1768 13144
rect 1820 13172 1826 13184
rect 2056 13181 2084 13280
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 4430 13308 4436 13320
rect 3467 13280 4436 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 4540 13317 4568 13348
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 4890 13376 4896 13388
rect 4847 13348 4896 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5258 13376 5264 13388
rect 5219 13348 5264 13376
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 6270 13376 6276 13388
rect 6231 13348 6276 13376
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6822 13376 6828 13388
rect 6503 13348 6828 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 8202 13336 8208 13388
rect 8260 13376 8266 13388
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 8260 13348 8309 13376
rect 8260 13336 8266 13348
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13308 4583 13311
rect 5626 13308 5632 13320
rect 4571 13280 5632 13308
rect 4571 13277 4583 13280
rect 4525 13271 4583 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 9968 13317 9996 13416
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11425 13447 11483 13453
rect 11425 13444 11437 13447
rect 11112 13416 11437 13444
rect 11112 13404 11118 13416
rect 11425 13413 11437 13416
rect 11471 13444 11483 13447
rect 11882 13444 11888 13456
rect 11471 13416 11888 13444
rect 11471 13413 11483 13416
rect 11425 13407 11483 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 10873 13379 10931 13385
rect 10873 13345 10885 13379
rect 10919 13345 10931 13379
rect 11698 13376 11704 13388
rect 11659 13348 11704 13376
rect 10873 13339 10931 13345
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13308 10011 13311
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 9999 13280 10609 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 10597 13277 10609 13280
rect 10643 13277 10655 13311
rect 10888 13308 10916 13339
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13376 12771 13379
rect 17862 13376 17868 13388
rect 12759 13348 17868 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 19702 13308 19708 13320
rect 10888 13280 19708 13308
rect 10597 13271 10655 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 3326 13240 3332 13252
rect 2332 13212 3332 13240
rect 2332 13184 2360 13212
rect 3326 13200 3332 13212
rect 3384 13200 3390 13252
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6181 13243 6239 13249
rect 6181 13240 6193 13243
rect 5408 13212 6193 13240
rect 5408 13200 5414 13212
rect 6181 13209 6193 13212
rect 6227 13209 6239 13243
rect 6181 13203 6239 13209
rect 8205 13243 8263 13249
rect 8205 13209 8217 13243
rect 8251 13240 8263 13243
rect 8251 13212 10272 13240
rect 8251 13209 8263 13212
rect 8205 13203 8263 13209
rect 2041 13175 2099 13181
rect 2041 13172 2053 13175
rect 1820 13144 2053 13172
rect 1820 13132 1826 13144
rect 2041 13141 2053 13144
rect 2087 13141 2099 13175
rect 2041 13135 2099 13141
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 2314 13172 2320 13184
rect 2179 13144 2320 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2406 13132 2412 13184
rect 2464 13172 2470 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 2464 13144 2513 13172
rect 2464 13132 2470 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 2501 13135 2559 13141
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 4982 13172 4988 13184
rect 4663 13144 4988 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5500 13144 5825 13172
rect 5500 13132 5506 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 6914 13172 6920 13184
rect 6875 13144 6920 13172
rect 5813 13135 5871 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 10244 13181 10272 13212
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 12437 13243 12495 13249
rect 12437 13240 12449 13243
rect 11756 13212 12449 13240
rect 11756 13200 11762 13212
rect 12437 13209 12449 13212
rect 12483 13209 12495 13243
rect 12437 13203 12495 13209
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13141 10287 13175
rect 10229 13135 10287 13141
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 10744 13144 10789 13172
rect 10744 13132 10750 13144
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 13078 13172 13084 13184
rect 12584 13144 12629 13172
rect 13039 13144 13084 13172
rect 12584 13132 12590 13144
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 20901 13175 20959 13181
rect 20901 13172 20913 13175
rect 20772 13144 20913 13172
rect 20772 13132 20778 13144
rect 20901 13141 20913 13144
rect 20947 13141 20959 13175
rect 20901 13135 20959 13141
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 1949 12971 2007 12977
rect 1949 12968 1961 12971
rect 1728 12940 1961 12968
rect 1728 12928 1734 12940
rect 1949 12937 1961 12940
rect 1995 12937 2007 12971
rect 1949 12931 2007 12937
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12937 2467 12971
rect 2409 12931 2467 12937
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12937 3111 12971
rect 3053 12931 3111 12937
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12968 5687 12971
rect 7377 12971 7435 12977
rect 7377 12968 7389 12971
rect 5675 12940 7389 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 7377 12937 7389 12940
rect 7423 12937 7435 12971
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7377 12931 7435 12937
rect 2424 12900 2452 12931
rect 2866 12900 2872 12912
rect 1688 12872 2452 12900
rect 2516 12872 2872 12900
rect 1688 12841 1716 12872
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2516 12832 2544 12872
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 2179 12804 2544 12832
rect 2593 12835 2651 12841
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 3068 12832 3096 12931
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 11054 12968 11060 12980
rect 8527 12940 11060 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 6880 12872 7972 12900
rect 6880 12860 6886 12872
rect 2639 12804 3096 12832
rect 3237 12835 3295 12841
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 4338 12832 4344 12844
rect 3283 12804 4344 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 5718 12764 5724 12776
rect 5679 12736 5724 12764
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12733 5871 12767
rect 6638 12764 6644 12776
rect 6599 12736 6644 12764
rect 5813 12727 5871 12733
rect 14 12656 20 12708
rect 72 12696 78 12708
rect 3881 12699 3939 12705
rect 3881 12696 3893 12699
rect 72 12668 3893 12696
rect 72 12656 78 12668
rect 3881 12665 3893 12668
rect 3927 12665 3939 12699
rect 3881 12659 3939 12665
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 4948 12668 5396 12696
rect 4948 12656 4954 12668
rect 3326 12588 3332 12640
rect 3384 12628 3390 12640
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 3384 12600 3525 12628
rect 3384 12588 3390 12600
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 4798 12588 4804 12640
rect 4856 12628 4862 12640
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 4856 12600 5273 12628
rect 4856 12588 4862 12600
rect 5261 12597 5273 12600
rect 5307 12597 5319 12631
rect 5368 12628 5396 12668
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 5828 12696 5856 12727
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 7098 12764 7104 12776
rect 7059 12736 7104 12764
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 5684 12668 5856 12696
rect 5684 12656 5690 12668
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 7760 12696 7788 12795
rect 7944 12773 7972 12872
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8018 12764 8024 12776
rect 7975 12736 8024 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8202 12696 8208 12708
rect 6972 12668 8208 12696
rect 6972 12656 6978 12668
rect 8202 12656 8208 12668
rect 8260 12696 8266 12708
rect 8496 12696 8524 12931
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 12158 12968 12164 12980
rect 12119 12940 12164 12968
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12529 12971 12587 12977
rect 12529 12937 12541 12971
rect 12575 12968 12587 12971
rect 13078 12968 13084 12980
rect 12575 12940 13084 12968
rect 12575 12937 12587 12940
rect 12529 12931 12587 12937
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 12066 12900 12072 12912
rect 8260 12668 8524 12696
rect 8588 12872 12072 12900
rect 8260 12656 8266 12668
rect 8588 12628 8616 12872
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9122 12832 9128 12844
rect 9079 12804 9128 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9122 12792 9128 12804
rect 9180 12832 9186 12844
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 9180 12804 10149 12832
rect 9180 12792 9186 12804
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 9674 12764 9680 12776
rect 9539 12736 9680 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 10410 12764 10416 12776
rect 10091 12736 10416 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 5368 12600 8616 12628
rect 9968 12628 9996 12727
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12406 12736 12633 12764
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 12406 12696 12434 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 16758 12764 16764 12776
rect 12851 12736 16764 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 10551 12668 12434 12696
rect 20441 12699 20499 12705
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 20441 12665 20453 12699
rect 20487 12696 20499 12699
rect 21542 12696 21548 12708
rect 20487 12668 21548 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 18414 12628 18420 12640
rect 9968 12600 18420 12628
rect 5261 12591 5319 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 20714 12628 20720 12640
rect 20675 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12628 20778 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 20772 12600 21189 12628
rect 20772 12588 20778 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 21177 12591 21235 12597
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 5813 12427 5871 12433
rect 5813 12424 5825 12427
rect 5776 12396 5825 12424
rect 5776 12384 5782 12396
rect 5813 12393 5825 12396
rect 5859 12393 5871 12427
rect 5813 12387 5871 12393
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 6604 12396 6837 12424
rect 6604 12384 6610 12396
rect 6825 12393 6837 12396
rect 6871 12393 6883 12427
rect 8018 12424 8024 12436
rect 6825 12387 6883 12393
rect 7392 12396 8024 12424
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12356 1639 12359
rect 2498 12356 2504 12368
rect 1627 12328 2504 12356
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 2498 12316 2504 12328
rect 2556 12316 2562 12368
rect 7392 12356 7420 12396
rect 8018 12384 8024 12396
rect 8076 12384 8082 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 8536 12396 9321 12424
rect 8536 12384 8542 12396
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 9309 12387 9367 12393
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 13170 12424 13176 12436
rect 11848 12396 13176 12424
rect 11848 12384 11854 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 19058 12424 19064 12436
rect 13872 12396 19064 12424
rect 13872 12384 13878 12396
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 9950 12356 9956 12368
rect 3804 12328 6408 12356
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2685 12291 2743 12297
rect 2685 12288 2697 12291
rect 2648 12260 2697 12288
rect 2648 12248 2654 12260
rect 2685 12257 2697 12260
rect 2731 12257 2743 12291
rect 2685 12251 2743 12257
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 3694 12288 3700 12300
rect 2832 12260 3700 12288
rect 2832 12248 2838 12260
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2866 12220 2872 12232
rect 2547 12192 2872 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3326 12220 3332 12232
rect 3287 12192 3332 12220
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 2593 12155 2651 12161
rect 2593 12121 2605 12155
rect 2639 12152 2651 12155
rect 2774 12152 2780 12164
rect 2639 12124 2780 12152
rect 2639 12121 2651 12124
rect 2593 12115 2651 12121
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 2884 12152 2912 12180
rect 3804 12161 3832 12328
rect 4798 12288 4804 12300
rect 4759 12260 4804 12288
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 2884 12124 3801 12152
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 5000 12152 5028 12251
rect 6380 12220 6408 12328
rect 6472 12328 7420 12356
rect 7484 12328 9956 12356
rect 6472 12297 6500 12328
rect 7484 12297 7512 12328
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 8168 12260 8401 12288
rect 8168 12248 8174 12260
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9640 12260 9873 12288
rect 9640 12248 9646 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12288 11023 12291
rect 11054 12288 11060 12300
rect 11011 12260 11060 12288
rect 11011 12257 11023 12260
rect 10965 12251 11023 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 6914 12220 6920 12232
rect 6380 12192 6920 12220
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 7156 12192 7205 12220
rect 7156 12180 7162 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 8202 12220 8208 12232
rect 8163 12192 8208 12220
rect 7193 12183 7251 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 11698 12220 11704 12232
rect 9784 12192 11704 12220
rect 7742 12152 7748 12164
rect 5000 12124 7748 12152
rect 3789 12115 3847 12121
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 8018 12112 8024 12164
rect 8076 12152 8082 12164
rect 9784 12152 9812 12192
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 11839 12192 13461 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 12268 12164 12296 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 20530 12220 20536 12232
rect 17083 12192 17448 12220
rect 20491 12192 20536 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 8076 12124 9812 12152
rect 8076 12112 8082 12124
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 12038 12155 12096 12161
rect 12038 12152 12050 12155
rect 9916 12124 12050 12152
rect 9916 12112 9922 12124
rect 12038 12121 12050 12124
rect 12084 12121 12096 12155
rect 12038 12115 12096 12121
rect 12250 12112 12256 12164
rect 12308 12112 12314 12164
rect 14366 12152 14372 12164
rect 12406 12124 14372 12152
rect 2130 12084 2136 12096
rect 2091 12056 2136 12084
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 2740 12056 3157 12084
rect 2740 12044 2746 12056
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3145 12047 3203 12053
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 4982 12084 4988 12096
rect 4755 12056 4988 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5350 12084 5356 12096
rect 5311 12056 5356 12084
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 5902 12084 5908 12096
rect 5592 12056 5908 12084
rect 5592 12044 5598 12056
rect 5902 12044 5908 12056
rect 5960 12084 5966 12096
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 5960 12056 6193 12084
rect 5960 12044 5966 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 6273 12087 6331 12093
rect 6273 12053 6285 12087
rect 6319 12084 6331 12087
rect 6546 12084 6552 12096
rect 6319 12056 6552 12084
rect 6319 12053 6331 12056
rect 6273 12047 6331 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7432 12056 7849 12084
rect 7432 12044 7438 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 7837 12047 7895 12053
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 7984 12056 8309 12084
rect 7984 12044 7990 12056
rect 8297 12053 8309 12056
rect 8343 12053 8355 12087
rect 8297 12047 8355 12053
rect 9033 12087 9091 12093
rect 9033 12053 9045 12087
rect 9079 12084 9091 12087
rect 9122 12084 9128 12096
rect 9079 12056 9128 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9769 12087 9827 12093
rect 9769 12053 9781 12087
rect 9815 12084 9827 12087
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 9815 12056 10333 12084
rect 9815 12053 9827 12056
rect 9769 12047 9827 12053
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 10321 12047 10379 12053
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10652 12056 10701 12084
rect 10652 12044 10658 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 10836 12056 10881 12084
rect 10836 12044 10842 12056
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 12406 12084 12434 12124
rect 14366 12112 14372 12124
rect 14424 12112 14430 12164
rect 16758 12152 16764 12164
rect 16816 12161 16822 12164
rect 16816 12155 16850 12161
rect 16702 12124 16764 12152
rect 16758 12112 16764 12124
rect 16838 12152 16850 12155
rect 17310 12152 17316 12164
rect 16838 12124 17316 12152
rect 16838 12121 16850 12124
rect 16816 12115 16850 12121
rect 16816 12112 16822 12115
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 13170 12084 13176 12096
rect 12216 12056 12434 12084
rect 13083 12056 13176 12084
rect 12216 12044 12222 12056
rect 13170 12044 13176 12056
rect 13228 12084 13234 12096
rect 14274 12084 14280 12096
rect 13228 12056 14280 12084
rect 13228 12044 13234 12056
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 15654 12084 15660 12096
rect 15615 12056 15660 12084
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 17420 12093 17448 12192
rect 20530 12180 20536 12192
rect 20588 12220 20594 12232
rect 21450 12220 21456 12232
rect 20588 12192 21456 12220
rect 20588 12180 20594 12192
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 19889 12155 19947 12161
rect 19889 12121 19901 12155
rect 19935 12152 19947 12155
rect 20257 12155 20315 12161
rect 20257 12152 20269 12155
rect 19935 12124 20269 12152
rect 19935 12121 19947 12124
rect 19889 12115 19947 12121
rect 20257 12121 20269 12124
rect 20303 12152 20315 12155
rect 20714 12152 20720 12164
rect 20303 12124 20720 12152
rect 20303 12121 20315 12124
rect 20257 12115 20315 12121
rect 20714 12112 20720 12124
rect 20772 12152 20778 12164
rect 20772 12124 21404 12152
rect 20772 12112 20778 12124
rect 21376 12096 21404 12124
rect 17405 12087 17463 12093
rect 17405 12053 17417 12087
rect 17451 12084 17463 12087
rect 18322 12084 18328 12096
rect 17451 12056 18328 12084
rect 17451 12053 17463 12056
rect 17405 12047 17463 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 20993 12087 21051 12093
rect 20993 12053 21005 12087
rect 21039 12084 21051 12087
rect 21082 12084 21088 12096
rect 21039 12056 21088 12084
rect 21039 12053 21051 12056
rect 20993 12047 21051 12053
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 21358 12084 21364 12096
rect 21319 12056 21364 12084
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 2188 11852 2513 11880
rect 2188 11840 2194 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 2501 11843 2559 11849
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 3016 11852 3157 11880
rect 3016 11840 3022 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 4982 11880 4988 11892
rect 4943 11852 4988 11880
rect 3145 11843 3203 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5442 11880 5448 11892
rect 5403 11852 5448 11880
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6052 11852 6377 11880
rect 6052 11840 6058 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6638 11840 6644 11892
rect 6696 11880 6702 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 6696 11852 6745 11880
rect 6696 11840 6702 11852
rect 6733 11849 6745 11852
rect 6779 11849 6791 11883
rect 6733 11843 6791 11849
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 7374 11880 7380 11892
rect 6871 11852 7380 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7524 11852 7757 11880
rect 7524 11840 7530 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 7745 11843 7803 11849
rect 8205 11883 8263 11889
rect 8205 11849 8217 11883
rect 8251 11880 8263 11883
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8251 11852 8769 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 9214 11880 9220 11892
rect 9175 11852 9220 11880
rect 8757 11843 8815 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 9858 11880 9864 11892
rect 9815 11852 9864 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 2590 11772 2596 11824
rect 2648 11812 2654 11824
rect 4341 11815 4399 11821
rect 2648 11784 4292 11812
rect 2648 11772 2654 11784
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11744 1455 11747
rect 1486 11744 1492 11756
rect 1443 11716 1492 11744
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1486 11704 1492 11716
rect 1544 11744 1550 11756
rect 2958 11744 2964 11756
rect 1544 11716 2964 11744
rect 1544 11704 1550 11716
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3326 11744 3332 11756
rect 3287 11716 3332 11744
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 2590 11676 2596 11688
rect 2551 11648 2596 11676
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 2774 11685 2780 11688
rect 2731 11679 2780 11685
rect 2731 11645 2743 11679
rect 2777 11645 2780 11679
rect 2731 11639 2780 11645
rect 2774 11636 2780 11639
rect 2832 11636 2838 11688
rect 4264 11676 4292 11784
rect 4341 11781 4353 11815
rect 4387 11812 4399 11815
rect 5350 11812 5356 11824
rect 4387 11784 5212 11812
rect 5311 11784 5356 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11744 4491 11747
rect 4614 11744 4620 11756
rect 4479 11716 4620 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 5184 11744 5212 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 9784 11812 9812 11843
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 15562 11880 15568 11892
rect 10008 11852 13676 11880
rect 15523 11852 15568 11880
rect 10008 11840 10014 11852
rect 13354 11812 13360 11824
rect 9048 11784 9812 11812
rect 9876 11784 13360 11812
rect 5902 11744 5908 11756
rect 5184 11716 5908 11744
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8662 11744 8668 11756
rect 8159 11716 8668 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 4525 11679 4583 11685
rect 4525 11676 4537 11679
rect 4264 11648 4537 11676
rect 4525 11645 4537 11648
rect 4571 11645 4583 11679
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 4525 11639 4583 11645
rect 3786 11568 3792 11620
rect 3844 11608 3850 11620
rect 3973 11611 4031 11617
rect 3973 11608 3985 11611
rect 3844 11580 3985 11608
rect 3844 11568 3850 11580
rect 3973 11577 3985 11580
rect 4019 11577 4031 11611
rect 4540 11608 4568 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7098 11676 7104 11688
rect 7055 11648 7104 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 9048 11676 9076 11784
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9876 11744 9904 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 10893 11747 10951 11753
rect 10893 11744 10905 11747
rect 9180 11716 9225 11744
rect 9324 11716 9904 11744
rect 9968 11716 10905 11744
rect 9180 11704 9186 11716
rect 8435 11648 9076 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 9324 11608 9352 11716
rect 9401 11679 9459 11685
rect 9401 11645 9413 11679
rect 9447 11676 9459 11679
rect 9968 11676 9996 11716
rect 10893 11713 10905 11716
rect 10939 11744 10951 11747
rect 11238 11744 11244 11756
rect 10939 11716 11244 11744
rect 10939 11713 10951 11716
rect 10893 11707 10951 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11698 11704 11704 11756
rect 11756 11744 11762 11756
rect 12325 11747 12383 11753
rect 12325 11744 12337 11747
rect 11756 11716 12337 11744
rect 11756 11704 11762 11716
rect 12325 11713 12337 11716
rect 12371 11744 12383 11747
rect 13170 11744 13176 11756
rect 12371 11716 13176 11744
rect 12371 11713 12383 11716
rect 12325 11707 12383 11713
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 9447 11648 9996 11676
rect 11149 11679 11207 11685
rect 9447 11645 9459 11648
rect 9401 11639 9459 11645
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 12069 11679 12127 11685
rect 11195 11648 11652 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 4540 11580 9352 11608
rect 3973 11571 4031 11577
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 2096 11512 2145 11540
rect 2096 11500 2102 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 3694 11540 3700 11552
rect 3607 11512 3700 11540
rect 2133 11503 2191 11509
rect 3694 11500 3700 11512
rect 3752 11540 3758 11552
rect 4154 11540 4160 11552
rect 3752 11512 4160 11540
rect 3752 11500 3758 11512
rect 4154 11500 4160 11512
rect 4212 11540 4218 11552
rect 7834 11540 7840 11552
rect 4212 11512 7840 11540
rect 4212 11500 4218 11512
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 11624 11549 11652 11648
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 11609 11543 11667 11549
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 12084 11540 12112 11639
rect 13648 11608 13676 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 19024 11852 19993 11880
rect 19024 11840 19030 11852
rect 19981 11849 19993 11852
rect 20027 11849 20039 11883
rect 19981 11843 20039 11849
rect 18322 11812 18328 11824
rect 14200 11784 15976 11812
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 14200 11753 14228 11784
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13780 11716 13829 11744
rect 13780 11704 13786 11716
rect 13817 11713 13829 11716
rect 13863 11744 13875 11747
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13863 11716 14197 11744
rect 13863 11713 13875 11716
rect 13817 11707 13875 11713
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 15948 11753 15976 11784
rect 16684 11784 18328 11812
rect 16684 11753 16712 11784
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 20806 11772 20812 11824
rect 20864 11812 20870 11824
rect 21094 11815 21152 11821
rect 21094 11812 21106 11815
rect 20864 11784 21106 11812
rect 20864 11772 20870 11784
rect 21094 11781 21106 11784
rect 21140 11781 21152 11815
rect 21094 11775 21152 11781
rect 14441 11747 14499 11753
rect 14441 11744 14453 11747
rect 14332 11716 14453 11744
rect 14332 11704 14338 11716
rect 14441 11713 14453 11716
rect 14487 11713 14499 11747
rect 14441 11707 14499 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 15979 11716 16313 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16301 11713 16313 11716
rect 16347 11744 16359 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16347 11716 16681 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16925 11747 16983 11753
rect 16925 11744 16937 11747
rect 16669 11707 16727 11713
rect 16776 11716 16937 11744
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 16776 11676 16804 11716
rect 16925 11713 16937 11716
rect 16971 11713 16983 11747
rect 18230 11744 18236 11756
rect 16925 11707 16983 11713
rect 17696 11716 18236 11744
rect 16540 11648 16804 11676
rect 16540 11636 16546 11648
rect 13648 11580 14228 11608
rect 12250 11540 12256 11552
rect 11655 11512 12256 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 13446 11540 13452 11552
rect 13359 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11540 13510 11552
rect 13814 11540 13820 11552
rect 13504 11512 13820 11540
rect 13504 11500 13510 11512
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14200 11540 14228 11580
rect 17696 11540 17724 11716
rect 18230 11704 18236 11716
rect 18288 11744 18294 11756
rect 18581 11747 18639 11753
rect 18581 11744 18593 11747
rect 18288 11716 18593 11744
rect 18288 11704 18294 11716
rect 18581 11713 18593 11716
rect 18627 11713 18639 11747
rect 21358 11744 21364 11756
rect 21319 11716 21364 11744
rect 18581 11707 18639 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 18322 11676 18328 11688
rect 18283 11648 18328 11676
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 14200 11512 17724 11540
rect 18049 11543 18107 11549
rect 18049 11509 18061 11543
rect 18095 11540 18107 11543
rect 18138 11540 18144 11552
rect 18095 11512 18144 11540
rect 18095 11509 18107 11512
rect 18049 11503 18107 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 19705 11543 19763 11549
rect 19705 11509 19717 11543
rect 19751 11540 19763 11543
rect 19794 11540 19800 11552
rect 19751 11512 19800 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2547 11308 2774 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2746 11268 2774 11308
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 3016 11308 3249 11336
rect 3016 11296 3022 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 3237 11299 3295 11305
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4488 11308 4537 11336
rect 4488 11296 4494 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12158 11336 12164 11348
rect 12115 11308 12164 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 12268 11308 14473 11336
rect 3050 11268 3056 11280
rect 2746 11240 3056 11268
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 5537 11271 5595 11277
rect 5537 11268 5549 11271
rect 5000 11240 5549 11268
rect 1946 11200 1952 11212
rect 1907 11172 1952 11200
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2038 11160 2044 11212
rect 2096 11200 2102 11212
rect 2096 11172 2141 11200
rect 2096 11160 2102 11172
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 2774 11200 2780 11212
rect 2648 11172 2780 11200
rect 2648 11160 2654 11172
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 5000 11209 5028 11240
rect 5537 11237 5549 11240
rect 5583 11237 5595 11271
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 5537 11231 5595 11237
rect 5920 11240 7849 11268
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5810 11200 5816 11212
rect 5215 11172 5816 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 5920 11141 5948 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 8202 11228 8208 11280
rect 8260 11268 8266 11280
rect 10594 11268 10600 11280
rect 8260 11240 10600 11268
rect 8260 11228 8266 11240
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11200 6239 11203
rect 6638 11200 6644 11212
rect 6227 11172 6644 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8076 11172 8401 11200
rect 8076 11160 8082 11172
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8720 11172 8953 11200
rect 8720 11160 8726 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 2280 11104 4169 11132
rect 2280 11092 2286 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11101 5963 11135
rect 7469 11135 7527 11141
rect 7469 11132 7481 11135
rect 5905 11095 5963 11101
rect 6748 11104 7481 11132
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 3476 11036 3801 11064
rect 3476 11024 3482 11036
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3789 11027 3847 11033
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 6748 11064 6776 11104
rect 7469 11101 7481 11104
rect 7515 11132 7527 11135
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 7515 11104 8217 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 8205 11101 8217 11104
rect 8251 11132 8263 11135
rect 9122 11132 9128 11144
rect 8251 11104 9128 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10962 11141 10968 11144
rect 10956 11095 10968 11141
rect 11020 11132 11026 11144
rect 12268 11132 12296 11308
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 14461 11299 14519 11305
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 16482 11336 16488 11348
rect 15528 11308 16488 11336
rect 15528 11296 15534 11308
rect 16482 11296 16488 11308
rect 16540 11336 16546 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 16540 11308 17509 11336
rect 16540 11296 16546 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 19116 11308 19349 11336
rect 19116 11296 19122 11308
rect 19337 11305 19349 11308
rect 19383 11336 19395 11339
rect 20806 11336 20812 11348
rect 19383 11308 20812 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 20806 11296 20812 11308
rect 20864 11296 20870 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 21358 11336 21364 11348
rect 21131 11308 21364 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12710 11268 12716 11280
rect 12391 11240 12716 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 13722 11160 13728 11172
rect 13780 11200 13786 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13780 11172 14105 11200
rect 13780 11160 13786 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 21100 11200 21128 11299
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 20763 11172 21128 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 11020 11104 12296 11132
rect 10962 11092 10968 11095
rect 11020 11092 11026 11104
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13228 11104 15516 11132
rect 13228 11092 13234 11104
rect 4856 11036 6776 11064
rect 4856 11024 4862 11036
rect 7098 11024 7104 11076
rect 7156 11064 7162 11076
rect 12158 11064 12164 11076
rect 7156 11036 10824 11064
rect 7156 11024 7162 11036
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 4890 10996 4896 11008
rect 2832 10968 2877 10996
rect 4851 10968 4896 10996
rect 2832 10956 2838 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6546 10996 6552 11008
rect 6052 10968 6097 10996
rect 6507 10968 6552 10996
rect 6052 10956 6058 10968
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 8202 10996 8208 11008
rect 6972 10968 8208 10996
rect 6972 10956 6978 10968
rect 8202 10956 8208 10968
rect 8260 10996 8266 11008
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 8260 10968 8309 10996
rect 8260 10956 8266 10968
rect 8297 10965 8309 10968
rect 8343 10965 8355 10999
rect 10796 10996 10824 11036
rect 11072 11036 12164 11064
rect 11072 10996 11100 11036
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 13458 11067 13516 11073
rect 13458 11064 13470 11067
rect 13412 11036 13470 11064
rect 13412 11024 13418 11036
rect 13458 11033 13470 11036
rect 13504 11033 13516 11067
rect 15488 11064 15516 11104
rect 15562 11092 15568 11144
rect 15620 11141 15626 11144
rect 15620 11132 15632 11141
rect 15841 11135 15899 11141
rect 15620 11104 15665 11132
rect 15620 11095 15632 11104
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 15887 11104 16129 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 16117 11101 16129 11104
rect 16163 11132 16175 11135
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 16163 11104 17877 11132
rect 16163 11101 16175 11104
rect 16117 11095 16175 11101
rect 17865 11101 17877 11104
rect 17911 11132 17923 11135
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17911 11104 18245 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 18233 11101 18245 11104
rect 18279 11132 18291 11135
rect 18322 11132 18328 11144
rect 18279 11104 18328 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 15620 11092 15626 11095
rect 18322 11092 18328 11104
rect 18380 11132 18386 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18380 11104 18613 11132
rect 18380 11092 18386 11104
rect 18601 11101 18613 11104
rect 18647 11132 18659 11135
rect 20732 11132 20760 11163
rect 18647 11104 20760 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 16390 11073 16396 11076
rect 16384 11064 16396 11073
rect 15488 11036 16252 11064
rect 16351 11036 16396 11064
rect 13458 11027 13516 11033
rect 10796 10968 11100 10996
rect 16224 10996 16252 11036
rect 16384 11027 16396 11036
rect 16390 11024 16396 11027
rect 16448 11024 16454 11076
rect 17034 11064 17040 11076
rect 16500 11036 17040 11064
rect 16500 10996 16528 11036
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 18966 11024 18972 11076
rect 19024 11064 19030 11076
rect 20450 11067 20508 11073
rect 20450 11064 20462 11067
rect 19024 11036 20462 11064
rect 19024 11024 19030 11036
rect 20450 11033 20462 11036
rect 20496 11033 20508 11067
rect 20450 11027 20508 11033
rect 16224 10968 16528 10996
rect 8297 10959 8355 10965
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1486 10752 1492 10804
rect 1544 10752 1550 10804
rect 1949 10795 2007 10801
rect 1949 10761 1961 10795
rect 1995 10792 2007 10795
rect 2130 10792 2136 10804
rect 1995 10764 2136 10792
rect 1995 10761 2007 10764
rect 1949 10755 2007 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2406 10792 2412 10804
rect 2367 10764 2412 10792
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3200 10764 3249 10792
rect 3200 10752 3206 10764
rect 3237 10761 3249 10764
rect 3283 10792 3295 10795
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 3283 10764 3801 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3789 10761 3801 10764
rect 3835 10792 3847 10795
rect 3970 10792 3976 10804
rect 3835 10764 3976 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4890 10792 4896 10804
rect 4295 10764 4896 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 7193 10795 7251 10801
rect 7193 10792 7205 10795
rect 5491 10764 7205 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 7193 10761 7205 10764
rect 7239 10761 7251 10795
rect 11146 10792 11152 10804
rect 7193 10755 7251 10761
rect 7300 10764 11152 10792
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 1504 10656 1532 10752
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2774 10724 2780 10736
rect 2363 10696 2780 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 6638 10724 6644 10736
rect 3712 10696 6644 10724
rect 2038 10656 2044 10668
rect 1443 10628 2044 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2590 10588 2596 10600
rect 2551 10560 2596 10588
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3712 10597 3740 10696
rect 6638 10684 6644 10696
rect 6696 10724 6702 10736
rect 7300 10724 7328 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 15654 10792 15660 10804
rect 14384 10764 15660 10792
rect 8938 10724 8944 10736
rect 6696 10696 7328 10724
rect 8899 10696 8944 10724
rect 6696 10684 6702 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 14216 10727 14274 10733
rect 14216 10693 14228 10727
rect 14262 10724 14274 10727
rect 14384 10724 14412 10764
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 18288 10764 18337 10792
rect 18288 10752 18294 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 14262 10696 14412 10724
rect 14476 10696 16160 10724
rect 14262 10693 14274 10696
rect 14216 10687 14274 10693
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 3970 10656 3976 10668
rect 3927 10628 3976 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4120 10628 5089 10656
rect 4120 10616 4126 10628
rect 5077 10625 5089 10628
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 6914 10656 6920 10668
rect 5776 10628 6920 10656
rect 5776 10616 5782 10628
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7331 10628 7941 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9306 10656 9312 10668
rect 8895 10628 9312 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 12250 10656 12256 10668
rect 12211 10628 12256 10656
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 14476 10665 14504 10696
rect 14461 10659 14519 10665
rect 12406 10628 14412 10656
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10557 3755 10591
rect 3697 10551 3755 10557
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 5442 10588 5448 10600
rect 5031 10560 5448 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 4908 10520 4936 10551
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10588 7159 10591
rect 8757 10591 8815 10597
rect 7147 10560 8708 10588
rect 7147 10557 7159 10560
rect 7101 10551 7159 10557
rect 6914 10520 6920 10532
rect 4908 10492 6920 10520
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 2406 10452 2412 10464
rect 1627 10424 2412 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5408 10424 5733 10452
rect 5408 10412 5414 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 6457 10455 6515 10461
rect 6457 10421 6469 10455
rect 6503 10452 6515 10455
rect 6822 10452 6828 10464
rect 6503 10424 6828 10452
rect 6503 10421 6515 10424
rect 6457 10415 6515 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7653 10455 7711 10461
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 8294 10452 8300 10464
rect 7699 10424 8300 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8680 10452 8708 10560
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 12406 10588 12434 10628
rect 8757 10551 8815 10557
rect 9140 10560 12434 10588
rect 14384 10588 14412 10628
rect 14461 10625 14473 10659
rect 14507 10625 14519 10659
rect 15470 10656 15476 10668
rect 14461 10619 14519 10625
rect 15120 10628 15476 10656
rect 15120 10588 15148 10628
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15838 10656 15844 10668
rect 15896 10665 15902 10668
rect 15808 10628 15844 10656
rect 15838 10616 15844 10628
rect 15896 10619 15908 10665
rect 15896 10616 15902 10619
rect 16132 10597 16160 10696
rect 18064 10696 21404 10724
rect 17770 10616 17776 10668
rect 17828 10665 17834 10668
rect 18064 10665 18092 10696
rect 17828 10656 17840 10665
rect 18049 10659 18107 10665
rect 17828 10628 17873 10656
rect 17828 10619 17840 10628
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 19449 10659 19507 10665
rect 19449 10625 19461 10659
rect 19495 10656 19507 10659
rect 19610 10656 19616 10668
rect 19495 10628 19616 10656
rect 19495 10625 19507 10628
rect 19449 10619 19507 10625
rect 17828 10616 17834 10619
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 19720 10665 19748 10696
rect 21376 10668 21404 10696
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 19794 10616 19800 10668
rect 19852 10656 19858 10668
rect 21094 10659 21152 10665
rect 21094 10656 21106 10659
rect 19852 10628 21106 10656
rect 19852 10616 19858 10628
rect 21094 10625 21106 10628
rect 21140 10625 21152 10659
rect 21358 10656 21364 10668
rect 21319 10628 21364 10656
rect 21094 10619 21152 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 14384 10560 15148 10588
rect 16117 10591 16175 10597
rect 8772 10520 8800 10551
rect 9140 10520 9168 10560
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16298 10588 16304 10600
rect 16163 10560 16304 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 8772 10492 9168 10520
rect 9232 10492 13584 10520
rect 9232 10452 9260 10492
rect 8680 10424 9260 10452
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9858 10452 9864 10464
rect 9355 10424 9864 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 12986 10452 12992 10464
rect 10284 10424 12992 10452
rect 10284 10412 10290 10424
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13446 10452 13452 10464
rect 13136 10424 13452 10452
rect 13136 10412 13142 10424
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 13556 10452 13584 10492
rect 14568 10492 15148 10520
rect 14568 10452 14596 10492
rect 14734 10452 14740 10464
rect 13556 10424 14596 10452
rect 14695 10424 14740 10452
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 15120 10452 15148 10492
rect 16390 10452 16396 10464
rect 15120 10424 16396 10452
rect 16390 10412 16396 10424
rect 16448 10452 16454 10464
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16448 10424 16681 10452
rect 16448 10412 16454 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 16669 10415 16727 10421
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19978 10452 19984 10464
rect 19116 10424 19984 10452
rect 19116 10412 19122 10424
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 1670 10248 1676 10260
rect 1627 10220 1676 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 4062 10248 4068 10260
rect 2087 10220 4068 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 6052 10220 6193 10248
rect 6052 10208 6058 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 7340 10220 8953 10248
rect 7340 10208 7346 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 11882 10248 11888 10260
rect 8941 10211 8999 10217
rect 10060 10220 11888 10248
rect 2130 10140 2136 10192
rect 2188 10180 2194 10192
rect 2314 10180 2320 10192
rect 2188 10152 2320 10180
rect 2188 10140 2194 10152
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 4154 10180 4160 10192
rect 3568 10152 4160 10180
rect 3568 10140 3574 10152
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 5810 10140 5816 10192
rect 5868 10180 5874 10192
rect 10060 10180 10088 10220
rect 11882 10208 11888 10220
rect 11940 10248 11946 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 11940 10220 12173 10248
rect 11940 10208 11946 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 17310 10248 17316 10260
rect 17271 10220 17316 10248
rect 12161 10211 12219 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 19058 10248 19064 10260
rect 17788 10220 19064 10248
rect 5868 10152 10088 10180
rect 5868 10140 5874 10152
rect 12986 10140 12992 10192
rect 13044 10180 13050 10192
rect 17788 10180 17816 10220
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 20993 10251 21051 10257
rect 20993 10248 21005 10251
rect 19260 10220 21005 10248
rect 13044 10152 17816 10180
rect 13044 10140 13050 10152
rect 3970 10112 3976 10124
rect 3931 10084 3976 10112
rect 3970 10072 3976 10084
rect 4028 10072 4034 10124
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5166 10112 5172 10124
rect 5123 10084 5172 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 8018 10112 8024 10124
rect 5675 10084 8024 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8389 10115 8447 10121
rect 8389 10112 8401 10115
rect 8260 10084 8401 10112
rect 8260 10072 8266 10084
rect 8389 10081 8401 10084
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9674 10112 9680 10124
rect 9631 10084 9680 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 19260 10121 19288 10220
rect 20993 10217 21005 10220
rect 21039 10248 21051 10251
rect 21358 10248 21364 10260
rect 21039 10220 21364 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 20625 10183 20683 10189
rect 20625 10149 20637 10183
rect 20671 10180 20683 10183
rect 20714 10180 20720 10192
rect 20671 10152 20720 10180
rect 20671 10149 20683 10152
rect 20625 10143 20683 10149
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 18693 10115 18751 10121
rect 18693 10081 18705 10115
rect 18739 10112 18751 10115
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 18739 10084 19257 10112
rect 18739 10081 18751 10084
rect 18693 10075 18751 10081
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 1360 10016 1409 10044
rect 1360 10004 1366 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1412 9976 1440 10007
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 1857 10047 1915 10053
rect 1857 10044 1869 10047
rect 1544 10016 1869 10044
rect 1544 10004 1550 10016
rect 1857 10013 1869 10016
rect 1903 10013 1915 10047
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 1857 10007 1915 10013
rect 2314 10004 2320 10016
rect 2372 10044 2378 10056
rect 2777 10047 2835 10053
rect 2777 10044 2789 10047
rect 2372 10016 2789 10044
rect 2372 10004 2378 10016
rect 2777 10013 2789 10016
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4120 10016 4905 10044
rect 4120 10004 4126 10016
rect 4893 10013 4905 10016
rect 4939 10044 4951 10047
rect 5718 10044 5724 10056
rect 4939 10016 5724 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 5828 10016 9321 10044
rect 1946 9976 1952 9988
rect 1412 9948 1952 9976
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 4798 9976 4804 9988
rect 3344 9948 4804 9976
rect 2498 9908 2504 9920
rect 2459 9880 2504 9908
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3344 9917 3372 9948
rect 4798 9936 4804 9948
rect 4856 9936 4862 9988
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 5828 9985 5856 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 10744 10016 10793 10044
rect 10744 10004 10750 10016
rect 10781 10013 10793 10016
rect 10827 10044 10839 10047
rect 12250 10044 12256 10056
rect 10827 10016 12256 10044
rect 10827 10013 10839 10016
rect 10781 10007 10839 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 18414 10004 18420 10056
rect 18472 10053 18478 10056
rect 18472 10044 18484 10053
rect 18472 10016 19748 10044
rect 18472 10007 18484 10016
rect 18472 10004 18478 10007
rect 19720 9988 19748 10016
rect 5813 9979 5871 9985
rect 5813 9976 5825 9979
rect 5592 9948 5825 9976
rect 5592 9936 5598 9948
rect 5813 9945 5825 9948
rect 5859 9945 5871 9979
rect 5813 9939 5871 9945
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 8297 9979 8355 9985
rect 8297 9976 8309 9979
rect 7156 9948 8309 9976
rect 7156 9936 7162 9948
rect 8297 9945 8309 9948
rect 8343 9945 8355 9979
rect 8297 9939 8355 9945
rect 11048 9979 11106 9985
rect 11048 9945 11060 9979
rect 11094 9976 11106 9979
rect 11146 9976 11152 9988
rect 11094 9948 11152 9976
rect 11094 9945 11106 9948
rect 11048 9939 11106 9945
rect 11146 9936 11152 9948
rect 11204 9976 11210 9988
rect 11698 9976 11704 9988
rect 11204 9948 11704 9976
rect 11204 9936 11210 9948
rect 11698 9936 11704 9948
rect 11756 9936 11762 9988
rect 16666 9976 16672 9988
rect 16579 9948 16672 9976
rect 16666 9936 16672 9948
rect 16724 9976 16730 9988
rect 19242 9976 19248 9988
rect 16724 9948 19248 9976
rect 16724 9936 16730 9948
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19490 9979 19548 9985
rect 19490 9976 19502 9979
rect 19392 9948 19502 9976
rect 19392 9936 19398 9948
rect 19490 9945 19502 9948
rect 19536 9945 19548 9979
rect 19490 9939 19548 9945
rect 19702 9936 19708 9988
rect 19760 9936 19766 9988
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 3108 9880 3341 9908
rect 3108 9868 3114 9880
rect 3329 9877 3341 9880
rect 3375 9877 3387 9911
rect 4430 9908 4436 9920
rect 4391 9880 4436 9908
rect 3329 9871 3387 9877
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4982 9868 4988 9920
rect 5040 9908 5046 9920
rect 5721 9911 5779 9917
rect 5721 9908 5733 9911
rect 5040 9880 5733 9908
rect 5040 9868 5046 9880
rect 5721 9877 5733 9880
rect 5767 9877 5779 9911
rect 5721 9871 5779 9877
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 5960 9880 6469 9908
rect 5960 9868 5966 9880
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6457 9871 6515 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7558 9908 7564 9920
rect 7519 9880 7564 9908
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7708 9880 7849 9908
rect 7708 9868 7714 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 7984 9880 8217 9908
rect 7984 9868 7990 9880
rect 8205 9877 8217 9880
rect 8251 9908 8263 9911
rect 8386 9908 8392 9920
rect 8251 9880 8392 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 9950 9908 9956 9920
rect 9456 9880 9501 9908
rect 9911 9880 9956 9908
rect 9456 9868 9462 9880
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 12250 9868 12256 9920
rect 12308 9908 12314 9920
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12308 9880 12541 9908
rect 12308 9868 12314 9880
rect 12529 9877 12541 9880
rect 12575 9908 12587 9911
rect 12802 9908 12808 9920
rect 12575 9880 12808 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 14645 9911 14703 9917
rect 14645 9877 14657 9911
rect 14691 9908 14703 9911
rect 16298 9908 16304 9920
rect 14691 9880 16304 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 17037 9911 17095 9917
rect 17037 9877 17049 9911
rect 17083 9908 17095 9911
rect 20162 9908 20168 9920
rect 17083 9880 20168 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 2685 9707 2743 9713
rect 2685 9704 2697 9707
rect 1544 9676 2697 9704
rect 1544 9664 1550 9676
rect 2685 9673 2697 9676
rect 2731 9673 2743 9707
rect 2685 9667 2743 9673
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7616 9676 7757 9704
rect 7616 9664 7622 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 9950 9704 9956 9716
rect 9815 9676 9956 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 19334 9704 19340 9716
rect 11112 9676 19340 9704
rect 11112 9664 11118 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 20898 9704 20904 9716
rect 19444 9676 20904 9704
rect 2038 9596 2044 9648
rect 2096 9636 2102 9648
rect 2317 9639 2375 9645
rect 2317 9636 2329 9639
rect 2096 9608 2329 9636
rect 2096 9596 2102 9608
rect 2317 9605 2329 9608
rect 2363 9605 2375 9639
rect 2317 9599 2375 9605
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 3142 9636 3148 9648
rect 2556 9608 3148 9636
rect 2556 9596 2562 9608
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 5077 9639 5135 9645
rect 5077 9636 5089 9639
rect 4120 9608 5089 9636
rect 4120 9596 4126 9608
rect 5077 9605 5089 9608
rect 5123 9605 5135 9639
rect 5077 9599 5135 9605
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 6914 9636 6920 9648
rect 6779 9608 6920 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 8386 9636 8392 9648
rect 8347 9608 8392 9636
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 9858 9636 9864 9648
rect 9819 9608 9864 9636
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 12434 9636 12440 9648
rect 9968 9608 12440 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 1854 9568 1860 9580
rect 1815 9540 1860 9568
rect 1854 9528 1860 9540
rect 1912 9568 1918 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 1912 9540 3065 9568
rect 1912 9528 1918 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3292 9540 3893 9568
rect 3292 9528 3298 9540
rect 3881 9537 3893 9540
rect 3927 9537 3939 9571
rect 4982 9568 4988 9580
rect 4943 9540 4988 9568
rect 3881 9531 3939 9537
rect 4982 9528 4988 9540
rect 5040 9568 5046 9580
rect 5534 9568 5540 9580
rect 5040 9540 5540 9568
rect 5040 9528 5046 9540
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7650 9568 7656 9580
rect 6871 9540 7656 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 1412 9500 1440 9528
rect 2774 9500 2780 9512
rect 1412 9472 2780 9500
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3142 9500 3148 9512
rect 2924 9472 3148 9500
rect 2924 9460 2930 9472
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3970 9500 3976 9512
rect 3931 9472 3976 9500
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4154 9500 4160 9512
rect 4111 9472 4160 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 5166 9500 5172 9512
rect 5127 9472 5172 9500
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5552 9500 5580 9528
rect 6914 9500 6920 9512
rect 5552 9472 6776 9500
rect 6875 9472 6920 9500
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 1627 9404 2774 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 2038 9364 2044 9376
rect 1999 9336 2044 9364
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 2746 9364 2774 9404
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3513 9435 3571 9441
rect 3513 9432 3525 9435
rect 3384 9404 3525 9432
rect 3384 9392 3390 9404
rect 3513 9401 3525 9404
rect 3559 9401 3571 9435
rect 3513 9395 3571 9401
rect 5258 9392 5264 9444
rect 5316 9432 5322 9444
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 5316 9404 6377 9432
rect 5316 9392 5322 9404
rect 6365 9401 6377 9404
rect 6411 9401 6423 9435
rect 6365 9395 6423 9401
rect 4522 9364 4528 9376
rect 2746 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4706 9364 4712 9376
rect 4663 9336 4712 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 4982 9324 4988 9376
rect 5040 9364 5046 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5040 9336 5641 9364
rect 5040 9324 5046 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 6748 9364 6776 9472
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 9968 9509 9996 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 12652 9639 12710 9645
rect 12652 9636 12664 9639
rect 12544 9608 12664 9636
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10652 9540 10793 9568
rect 10652 9528 10658 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 12544 9568 12572 9608
rect 12652 9605 12664 9608
rect 12698 9636 12710 9639
rect 14734 9636 14740 9648
rect 12698 9608 14740 9636
rect 12698 9605 12710 9608
rect 12652 9599 12710 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 15562 9636 15568 9648
rect 15475 9608 15568 9636
rect 15562 9596 15568 9608
rect 15620 9636 15626 9648
rect 16298 9636 16304 9648
rect 15620 9608 16304 9636
rect 15620 9596 15626 9608
rect 16298 9596 16304 9608
rect 16356 9636 16362 9648
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16356 9608 16773 9636
rect 16356 9596 16362 9608
rect 16761 9605 16773 9608
rect 16807 9636 16819 9639
rect 16807 9608 18460 9636
rect 16807 9605 16819 9608
rect 16761 9599 16819 9605
rect 18432 9580 18460 9608
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 19444 9636 19472 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 21358 9704 21364 9716
rect 21319 9676 21364 9704
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 19300 9608 19472 9636
rect 19300 9596 19306 9608
rect 19978 9596 19984 9648
rect 20036 9636 20042 9648
rect 20450 9639 20508 9645
rect 20450 9636 20462 9639
rect 20036 9608 20462 9636
rect 20036 9596 20042 9608
rect 20450 9605 20462 9608
rect 20496 9605 20508 9639
rect 20450 9599 20508 9605
rect 12216 9540 12572 9568
rect 12216 9528 12222 9540
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12952 9540 13185 9568
rect 12952 9528 12958 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 18138 9528 18144 9580
rect 18196 9577 18202 9580
rect 18196 9568 18208 9577
rect 18414 9568 18420 9580
rect 18196 9540 18241 9568
rect 18327 9540 18420 9568
rect 18196 9531 18208 9540
rect 18196 9528 18202 9531
rect 18414 9528 18420 9540
rect 18472 9568 18478 9580
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 18472 9540 18889 9568
rect 18472 9528 18478 9540
rect 18877 9537 18889 9540
rect 18923 9568 18935 9571
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 18923 9540 20729 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 20717 9537 20729 9540
rect 20763 9568 20775 9571
rect 21376 9568 21404 9664
rect 20763 9540 21404 9568
rect 20763 9537 20775 9540
rect 20717 9531 20775 9537
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 9953 9503 10011 9509
rect 8067 9472 9674 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 7064 9404 7389 9432
rect 7064 9392 7070 9404
rect 7377 9401 7389 9404
rect 7423 9401 7435 9435
rect 7852 9432 7880 9463
rect 9646 9432 9674 9472
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 10870 9500 10876 9512
rect 9953 9463 10011 9469
rect 10336 9472 10741 9500
rect 10831 9472 10876 9500
rect 10336 9432 10364 9472
rect 7852 9404 9536 9432
rect 9646 9404 10364 9432
rect 10413 9435 10471 9441
rect 7377 9395 7435 9401
rect 7558 9364 7564 9376
rect 6748 9336 7564 9364
rect 5629 9327 5687 9333
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9180 9336 9413 9364
rect 9180 9324 9186 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9508 9364 9536 9404
rect 10413 9401 10425 9435
rect 10459 9401 10471 9435
rect 10713 9432 10741 9472
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 11054 9500 11060 9512
rect 11015 9472 11060 9500
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 10713 9404 12020 9432
rect 10413 9395 10471 9401
rect 10428 9364 10456 9395
rect 9508 9336 10456 9364
rect 9401 9327 9459 9333
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11296 9336 11529 9364
rect 11296 9324 11302 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11992 9364 12020 9404
rect 13170 9392 13176 9444
rect 13228 9432 13234 9444
rect 17034 9432 17040 9444
rect 13228 9404 16896 9432
rect 16995 9404 17040 9432
rect 13228 9392 13234 9404
rect 12618 9364 12624 9376
rect 11992 9336 12624 9364
rect 11517 9327 11575 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15804 9336 15853 9364
rect 15804 9324 15810 9336
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 16868 9364 16896 9404
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 19518 9364 19524 9376
rect 16868 9336 19524 9364
rect 15841 9327 15899 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4028 9132 4261 9160
rect 4028 9120 4034 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 4448 9132 6868 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 4448 9092 4476 9132
rect 6840 9092 6868 9132
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 6972 9132 11284 9160
rect 6972 9120 6978 9132
rect 7926 9092 7932 9104
rect 1627 9064 4476 9092
rect 4540 9064 4936 9092
rect 6840 9064 7932 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 4540 9024 4568 9064
rect 4706 9024 4712 9036
rect 2731 8996 4568 9024
rect 4667 8996 4712 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 4908 9033 4936 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7650 9024 7656 9036
rect 6963 8996 7656 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 2648 8928 3801 8956
rect 2648 8916 2654 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4488 8928 4629 8956
rect 4488 8916 4494 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4908 8956 4936 8987
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8067 8996 9812 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8662 8956 8668 8968
rect 4908 8928 8668 8956
rect 4617 8919 4675 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 1412 8888 1440 8916
rect 3326 8888 3332 8900
rect 1412 8860 3332 8888
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 5721 8891 5779 8897
rect 5721 8888 5733 8891
rect 4448 8860 5733 8888
rect 4448 8832 4476 8860
rect 5721 8857 5733 8860
rect 5767 8857 5779 8891
rect 5721 8851 5779 8857
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 6052 8860 6469 8888
rect 6052 8848 6058 8860
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 6788 8860 7849 8888
rect 6788 8848 6794 8860
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 7837 8851 7895 8857
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2498 8820 2504 8832
rect 2372 8792 2504 8820
rect 2372 8780 2378 8792
rect 2498 8780 2504 8792
rect 2556 8820 2562 8832
rect 2777 8823 2835 8829
rect 2777 8820 2789 8823
rect 2556 8792 2789 8820
rect 2556 8780 2562 8792
rect 2777 8789 2789 8792
rect 2823 8789 2835 8823
rect 2777 8783 2835 8789
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 2924 8792 2969 8820
rect 2924 8780 2930 8792
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 3973 8823 4031 8829
rect 3973 8820 3985 8823
rect 3936 8792 3985 8820
rect 3936 8780 3942 8792
rect 3973 8789 3985 8792
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 4430 8780 4436 8832
rect 4488 8780 4494 8832
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5684 8792 6101 8820
rect 5684 8780 5690 8792
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 6089 8783 6147 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 7745 8823 7803 8829
rect 7745 8820 7757 8823
rect 7616 8792 7757 8820
rect 7616 8780 7622 8792
rect 7745 8789 7757 8792
rect 7791 8789 7803 8823
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 7745 8783 7803 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8812 8792 8953 8820
rect 8812 8780 8818 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 9490 8820 9496 8832
rect 9451 8792 9496 8820
rect 8941 8783 8999 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9784 8829 9812 8996
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 10882 8959 10940 8965
rect 10882 8956 10894 8959
rect 10560 8928 10894 8956
rect 10560 8916 10566 8928
rect 10882 8925 10894 8928
rect 10928 8956 10940 8959
rect 11146 8956 11152 8968
rect 10928 8928 11008 8956
rect 11107 8928 11152 8956
rect 10928 8925 10940 8928
rect 10882 8919 10940 8925
rect 9769 8823 9827 8829
rect 9769 8789 9781 8823
rect 9815 8820 9827 8823
rect 10594 8820 10600 8832
rect 9815 8792 10600 8820
rect 9815 8789 9827 8792
rect 9769 8783 9827 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10980 8820 11008 8928
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11256 8956 11284 9132
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11790 9160 11796 9172
rect 11388 9132 11796 9160
rect 11388 9120 11394 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 15930 9160 15936 9172
rect 15891 9132 15936 9160
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 17681 9163 17739 9169
rect 17681 9129 17693 9163
rect 17727 9160 17739 9163
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 17727 9132 18245 9160
rect 17727 9129 17739 9132
rect 17681 9123 17739 9129
rect 18233 9129 18245 9132
rect 18279 9160 18291 9163
rect 18414 9160 18420 9172
rect 18279 9132 18420 9160
rect 18279 9129 18291 9132
rect 18233 9123 18291 9129
rect 15562 9024 15568 9036
rect 15523 8996 15568 9024
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 17313 9027 17371 9033
rect 17313 8993 17325 9027
rect 17359 9024 17371 9027
rect 17696 9024 17724 9123
rect 18414 9120 18420 9132
rect 18472 9160 18478 9172
rect 18509 9163 18567 9169
rect 18509 9160 18521 9163
rect 18472 9132 18521 9160
rect 18472 9120 18478 9132
rect 18509 9129 18521 9132
rect 18555 9160 18567 9163
rect 19337 9163 19395 9169
rect 19337 9160 19349 9163
rect 18555 9132 19349 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 19337 9129 19349 9132
rect 19383 9129 19395 9163
rect 19702 9160 19708 9172
rect 19663 9132 19708 9160
rect 19337 9123 19395 9129
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 17359 8996 17724 9024
rect 21085 9027 21143 9033
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 21085 8993 21097 9027
rect 21131 9024 21143 9027
rect 21358 9024 21364 9036
rect 21131 8996 21364 9024
rect 21131 8993 21143 8996
rect 21085 8987 21143 8993
rect 21358 8984 21364 8996
rect 21416 8984 21422 9036
rect 12802 8956 12808 8968
rect 11256 8928 12684 8956
rect 12763 8928 12808 8956
rect 12066 8848 12072 8900
rect 12124 8888 12130 8900
rect 12538 8891 12596 8897
rect 12538 8888 12550 8891
rect 12124 8860 12550 8888
rect 12124 8848 12130 8860
rect 12538 8857 12550 8860
rect 12584 8857 12596 8891
rect 12656 8888 12684 8928
rect 12802 8916 12808 8928
rect 12860 8956 12866 8968
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12860 8928 13093 8956
rect 12860 8916 12866 8928
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 15298 8959 15356 8965
rect 15298 8956 15310 8959
rect 13872 8928 15310 8956
rect 13872 8916 13878 8928
rect 15298 8925 15310 8928
rect 15344 8925 15356 8959
rect 15298 8919 15356 8925
rect 20806 8916 20812 8968
rect 20864 8965 20870 8968
rect 20864 8956 20876 8965
rect 20864 8928 20909 8956
rect 20864 8919 20876 8928
rect 20864 8916 20870 8919
rect 12986 8888 12992 8900
rect 12656 8860 12992 8888
rect 12538 8851 12596 8857
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 14642 8888 14648 8900
rect 14108 8860 14648 8888
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 10980 8792 11437 8820
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 14108 8820 14136 8860
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 17068 8891 17126 8897
rect 17068 8857 17080 8891
rect 17114 8888 17126 8891
rect 17954 8888 17960 8900
rect 17114 8860 17960 8888
rect 17114 8857 17126 8860
rect 17068 8851 17126 8857
rect 17954 8848 17960 8860
rect 18012 8848 18018 8900
rect 11848 8792 14136 8820
rect 14185 8823 14243 8829
rect 11848 8780 11854 8792
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 14274 8820 14280 8832
rect 14231 8792 14280 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 15746 8780 15752 8832
rect 15804 8820 15810 8832
rect 20622 8820 20628 8832
rect 15804 8792 20628 8820
rect 15804 8780 15810 8792
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5258 8616 5264 8628
rect 5219 8588 5264 8616
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 8386 8616 8392 8628
rect 7515 8588 8392 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8536 8588 9413 8616
rect 8536 8576 8542 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 9548 8588 9781 8616
rect 9548 8576 9554 8588
rect 9769 8585 9781 8588
rect 9815 8585 9827 8619
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 9769 8579 9827 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 13354 8616 13360 8628
rect 13315 8588 13360 8616
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 15105 8619 15163 8625
rect 13504 8588 13952 8616
rect 13504 8576 13510 8588
rect 1854 8508 1860 8560
rect 1912 8548 1918 8560
rect 3329 8551 3387 8557
rect 3329 8548 3341 8551
rect 1912 8520 3341 8548
rect 1912 8508 1918 8520
rect 3329 8517 3341 8520
rect 3375 8517 3387 8551
rect 3329 8511 3387 8517
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 3936 8520 4476 8548
rect 3936 8508 3942 8520
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 4246 8480 4252 8492
rect 4207 8452 4252 8480
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2314 8412 2320 8424
rect 1728 8384 2320 8412
rect 1728 8372 1734 8384
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 4338 8412 4344 8424
rect 2746 8384 4200 8412
rect 4299 8384 4344 8412
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2746 8344 2774 8384
rect 1627 8316 2774 8344
rect 3881 8347 3939 8353
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4062 8344 4068 8356
rect 3927 8316 4068 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4172 8344 4200 8384
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4448 8421 4476 8520
rect 4522 8508 4528 8560
rect 4580 8548 4586 8560
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 4580 8520 5365 8548
rect 4580 8508 4586 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 10962 8548 10968 8560
rect 5353 8511 5411 8517
rect 6748 8520 10968 8548
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 6748 8480 6776 8520
rect 10962 8508 10968 8520
rect 11020 8508 11026 8560
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 12814 8551 12872 8557
rect 12814 8548 12826 8551
rect 11940 8520 12826 8548
rect 11940 8508 11946 8520
rect 12814 8517 12826 8520
rect 12860 8517 12872 8551
rect 13170 8548 13176 8560
rect 12814 8511 12872 8517
rect 12912 8520 13176 8548
rect 5224 8452 6776 8480
rect 6825 8483 6883 8489
rect 5224 8440 5230 8452
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 6871 8452 8493 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 12912 8480 12940 8520
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 13924 8548 13952 8588
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15194 8616 15200 8628
rect 15151 8588 15200 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15194 8576 15200 8588
rect 15252 8616 15258 8628
rect 15562 8616 15568 8628
rect 15252 8588 15568 8616
rect 15252 8576 15258 8588
rect 15562 8576 15568 8588
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8616 15715 8619
rect 15930 8616 15936 8628
rect 15703 8588 15936 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 15930 8576 15936 8588
rect 15988 8616 15994 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 15988 8588 16221 8616
rect 15988 8576 15994 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 16209 8579 16267 8585
rect 13924 8520 15424 8548
rect 8720 8452 12940 8480
rect 8720 8440 8726 8452
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 13044 8452 13093 8480
rect 13044 8440 13050 8452
rect 13081 8449 13093 8452
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14470 8483 14528 8489
rect 14470 8480 14482 8483
rect 13780 8452 14482 8480
rect 13780 8440 13786 8452
rect 14470 8449 14482 8452
rect 14516 8480 14528 8483
rect 14737 8483 14795 8489
rect 14516 8452 14688 8480
rect 14516 8449 14528 8452
rect 14470 8443 14528 8449
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5626 8412 5632 8424
rect 5583 8384 5632 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8294 8412 8300 8424
rect 7791 8384 8300 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 9858 8412 9864 8424
rect 9819 8384 9864 8412
rect 8757 8375 8815 8381
rect 5718 8344 5724 8356
rect 4172 8316 5724 8344
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5868 8316 5917 8344
rect 5868 8304 5874 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 5905 8307 5963 8313
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 6972 8316 7113 8344
rect 6972 8304 6978 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 8772 8344 8800 8375
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 11882 8412 11888 8424
rect 10091 8384 11888 8412
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 14660 8412 14688 8452
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15194 8480 15200 8492
rect 14783 8452 15200 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 15286 8412 15292 8424
rect 14660 8384 15292 8412
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15396 8412 15424 8520
rect 16224 8480 16252 8579
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17920 8588 18061 8616
rect 17920 8576 17926 8588
rect 18049 8585 18061 8588
rect 18095 8616 18107 8619
rect 18095 8588 20116 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 17586 8548 17592 8560
rect 16684 8520 17592 8548
rect 16684 8489 16712 8520
rect 17586 8508 17592 8520
rect 17644 8548 17650 8560
rect 20088 8548 20116 8588
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21232 8588 21373 8616
rect 21232 8576 21238 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 20226 8551 20284 8557
rect 20226 8548 20238 8551
rect 17644 8520 20024 8548
rect 20088 8520 20238 8548
rect 17644 8508 17650 8520
rect 18340 8489 18368 8520
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16224 8452 16681 8480
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16925 8483 16983 8489
rect 16925 8480 16937 8483
rect 16669 8443 16727 8449
rect 16776 8452 16937 8480
rect 16776 8412 16804 8452
rect 16925 8449 16937 8452
rect 16971 8449 16983 8483
rect 16925 8443 16983 8449
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 19996 8489 20024 8520
rect 20226 8517 20238 8520
rect 20272 8517 20284 8551
rect 20226 8511 20284 8517
rect 18581 8483 18639 8489
rect 18581 8480 18593 8483
rect 18472 8452 18593 8480
rect 18472 8440 18478 8452
rect 18581 8449 18593 8452
rect 18627 8449 18639 8483
rect 18581 8443 18639 8449
rect 19981 8483 20039 8489
rect 19981 8449 19993 8483
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 15396 8384 16804 8412
rect 11790 8344 11796 8356
rect 8772 8316 11796 8344
rect 7101 8307 7159 8313
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 12066 8344 12072 8356
rect 11900 8316 12072 8344
rect 4890 8276 4896 8288
rect 4851 8248 4896 8276
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 8113 8279 8171 8285
rect 8113 8276 8125 8279
rect 7524 8248 8125 8276
rect 7524 8236 7530 8248
rect 8113 8245 8125 8248
rect 8159 8245 8171 8279
rect 8113 8239 8171 8245
rect 11701 8279 11759 8285
rect 11701 8245 11713 8279
rect 11747 8276 11759 8279
rect 11900 8276 11928 8316
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 19518 8304 19524 8356
rect 19576 8344 19582 8356
rect 19705 8347 19763 8353
rect 19705 8344 19717 8347
rect 19576 8316 19717 8344
rect 19576 8304 19582 8316
rect 19705 8313 19717 8316
rect 19751 8313 19763 8347
rect 19705 8307 19763 8313
rect 11747 8248 11928 8276
rect 11747 8245 11759 8248
rect 11701 8239 11759 8245
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 15838 8276 15844 8288
rect 12216 8248 15844 8276
rect 12216 8236 12222 8248
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 1452 8044 3801 8072
rect 1452 8032 1458 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4246 8072 4252 8084
rect 4203 8044 4252 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 4356 8044 6193 8072
rect 4356 8004 4384 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7558 8072 7564 8084
rect 7239 8044 7564 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 8570 8072 8576 8084
rect 7668 8044 8576 8072
rect 5905 8007 5963 8013
rect 1872 7976 4384 8004
rect 4448 7976 5672 8004
rect 1872 7880 1900 7976
rect 4448 7936 4476 7976
rect 1964 7908 4476 7936
rect 4801 7939 4859 7945
rect 1394 7828 1400 7880
rect 1452 7877 1458 7880
rect 1452 7871 1479 7877
rect 1467 7868 1479 7871
rect 1854 7868 1860 7880
rect 1467 7840 1716 7868
rect 1767 7840 1860 7868
rect 1467 7837 1479 7840
rect 1452 7831 1479 7837
rect 1452 7828 1458 7831
rect 1688 7800 1716 7840
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 1964 7800 1992 7908
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 5166 7936 5172 7948
rect 4847 7908 5172 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 5445 7939 5503 7945
rect 5316 7908 5361 7936
rect 5316 7896 5322 7908
rect 5445 7905 5457 7939
rect 5491 7936 5503 7939
rect 5534 7936 5540 7948
rect 5491 7908 5540 7936
rect 5491 7905 5503 7908
rect 5445 7899 5503 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 5644 7936 5672 7976
rect 5905 7973 5917 8007
rect 5951 8004 5963 8007
rect 7668 8004 7696 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 9916 8044 10057 8072
rect 9916 8032 9922 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 10045 8035 10103 8041
rect 14292 8044 15332 8072
rect 5951 7976 7696 8004
rect 5951 7973 5963 7976
rect 5905 7967 5963 7973
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 8352 7976 11008 8004
rect 8352 7964 8358 7976
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 5644 7908 6561 7936
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 6549 7899 6607 7905
rect 6656 7908 7665 7936
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2682 7868 2688 7880
rect 2363 7840 2688 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3237 7871 3295 7877
rect 2832 7840 2877 7868
rect 2832 7828 2838 7840
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3326 7868 3332 7880
rect 3283 7840 3332 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7864 4583 7871
rect 4706 7864 4712 7880
rect 4571 7837 4712 7864
rect 4525 7836 4712 7837
rect 4525 7831 4583 7836
rect 4706 7828 4712 7836
rect 4764 7868 4770 7880
rect 6656 7868 6684 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7834 7936 7840 7948
rect 7795 7908 7840 7936
rect 7653 7899 7711 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7936 9551 7939
rect 9539 7908 10916 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 4764 7840 6684 7868
rect 4764 7828 4770 7840
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7340 7840 7573 7868
rect 7340 7828 7346 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 7561 7831 7619 7837
rect 7668 7840 9597 7868
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 1688 7772 1992 7800
rect 2056 7772 5549 7800
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1762 7732 1768 7744
rect 1627 7704 1768 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 2056 7741 2084 7772
rect 5537 7769 5549 7772
rect 5583 7769 5595 7803
rect 5537 7763 5595 7769
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 7668 7800 7696 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9766 7868 9772 7880
rect 9723 7840 9772 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 6880 7772 7696 7800
rect 6880 7760 6886 7772
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 10888 7800 10916 7908
rect 10980 7868 11008 7976
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11698 7936 11704 7948
rect 11296 7908 11704 7936
rect 11296 7896 11302 7908
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 14292 7936 14320 8044
rect 15304 8004 15332 8044
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 15436 8044 15669 8072
rect 15436 8032 15442 8044
rect 15657 8041 15669 8044
rect 15703 8072 15715 8075
rect 17310 8072 17316 8084
rect 15703 8044 16988 8072
rect 17271 8044 17316 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 15838 8004 15844 8016
rect 15304 7976 15844 8004
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 15930 7936 15936 7948
rect 12656 7908 14320 7936
rect 15891 7908 15936 7936
rect 12656 7868 12684 7908
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 10980 7840 12684 7868
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 12802 7868 12808 7880
rect 12759 7840 12808 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 12802 7828 12808 7840
rect 12860 7868 12866 7880
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12860 7840 13277 7868
rect 12860 7828 12866 7840
rect 13265 7837 13277 7840
rect 13311 7868 13323 7871
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 13311 7840 13645 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 13633 7837 13645 7840
rect 13679 7868 13691 7871
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13679 7840 14289 7868
rect 13679 7837 13691 7840
rect 13633 7831 13691 7837
rect 14277 7837 14289 7840
rect 14323 7868 14335 7871
rect 15948 7868 15976 7896
rect 14323 7840 15976 7868
rect 16960 7868 16988 8044
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 17586 8072 17592 8084
rect 17547 8044 17592 8072
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 19610 8072 19616 8084
rect 17736 8044 19616 8072
rect 17736 8032 17742 8044
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 20622 8072 20628 8084
rect 20583 8044 20628 8072
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 20993 8075 21051 8081
rect 20993 8041 21005 8075
rect 21039 8072 21051 8075
rect 21358 8072 21364 8084
rect 21039 8044 21364 8072
rect 21039 8041 21051 8044
rect 20993 8035 21051 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 17604 7936 17632 8032
rect 18506 8004 18512 8016
rect 18467 7976 18512 8004
rect 18506 7964 18512 7976
rect 18564 7964 18570 8016
rect 20640 8004 20668 8032
rect 21266 8004 21272 8016
rect 20640 7976 21272 8004
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 17604 7908 19257 7936
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 16960 7840 18153 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 18141 7837 18153 7840
rect 18187 7868 18199 7871
rect 18414 7868 18420 7880
rect 18187 7840 18420 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 12468 7803 12526 7809
rect 8168 7772 10824 7800
rect 10888 7772 12434 7800
rect 8168 7760 8174 7772
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7701 2099 7735
rect 2041 7695 2099 7701
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 2958 7732 2964 7744
rect 2547 7704 2964 7732
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4617 7735 4675 7741
rect 4617 7732 4629 7735
rect 4028 7704 4629 7732
rect 4028 7692 4034 7704
rect 4617 7701 4629 7704
rect 4663 7701 4675 7735
rect 8202 7732 8208 7744
rect 8163 7704 8208 7732
rect 4617 7695 4675 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8938 7732 8944 7744
rect 8899 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10686 7732 10692 7744
rect 10647 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 10796 7732 10824 7772
rect 11333 7735 11391 7741
rect 11333 7732 11345 7735
rect 10796 7704 11345 7732
rect 11333 7701 11345 7704
rect 11379 7732 11391 7735
rect 12158 7732 12164 7744
rect 11379 7704 12164 7732
rect 11379 7701 11391 7704
rect 11333 7695 11391 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12406 7732 12434 7772
rect 12468 7769 12480 7803
rect 12514 7800 12526 7803
rect 12618 7800 12624 7812
rect 12514 7772 12624 7800
rect 12514 7769 12526 7772
rect 12468 7763 12526 7769
rect 12618 7760 12624 7772
rect 12676 7800 12682 7812
rect 12894 7800 12900 7812
rect 12676 7772 12900 7800
rect 12676 7760 12682 7772
rect 12894 7760 12900 7772
rect 12952 7760 12958 7812
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 14522 7803 14580 7809
rect 14522 7800 14534 7803
rect 14424 7772 14534 7800
rect 14424 7760 14430 7772
rect 14522 7769 14534 7772
rect 14568 7769 14580 7803
rect 16200 7803 16258 7809
rect 16200 7800 16212 7803
rect 14522 7763 14580 7769
rect 15396 7772 16212 7800
rect 15396 7732 15424 7772
rect 16200 7769 16212 7772
rect 16246 7800 16258 7803
rect 16298 7800 16304 7812
rect 16246 7772 16304 7800
rect 16246 7769 16258 7772
rect 16200 7763 16258 7769
rect 16298 7760 16304 7772
rect 16356 7760 16362 7812
rect 19512 7803 19570 7809
rect 19512 7769 19524 7803
rect 19558 7800 19570 7803
rect 19610 7800 19616 7812
rect 19558 7772 19616 7800
rect 19558 7769 19570 7772
rect 19512 7763 19570 7769
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 12406 7704 15424 7732
rect 15838 7692 15844 7744
rect 15896 7732 15902 7744
rect 19702 7732 19708 7744
rect 15896 7704 19708 7732
rect 15896 7692 15902 7704
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 2498 7528 2504 7540
rect 2459 7500 2504 7528
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 2648 7500 3985 7528
rect 2648 7488 2654 7500
rect 3973 7497 3985 7500
rect 4019 7528 4031 7531
rect 4246 7528 4252 7540
rect 4019 7500 4252 7528
rect 4019 7497 4031 7500
rect 3973 7491 4031 7497
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4396 7500 4445 7528
rect 4396 7488 4402 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4948 7500 5089 7528
rect 4948 7488 4954 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5534 7528 5540 7540
rect 5316 7500 5540 7528
rect 5316 7488 5322 7500
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 7190 7528 7196 7540
rect 7147 7500 7196 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 8202 7528 8208 7540
rect 7515 7500 8208 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 10686 7528 10692 7540
rect 8312 7500 10692 7528
rect 4982 7460 4988 7472
rect 1412 7432 4988 7460
rect 1412 7404 1440 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 6733 7463 6791 7469
rect 6733 7460 6745 7463
rect 5500 7432 6745 7460
rect 5500 7420 5506 7432
rect 6733 7429 6745 7432
rect 6779 7429 6791 7463
rect 6733 7423 6791 7429
rect 7374 7420 7380 7472
rect 7432 7460 7438 7472
rect 7561 7463 7619 7469
rect 7561 7460 7573 7463
rect 7432 7432 7573 7460
rect 7432 7420 7438 7432
rect 7561 7429 7573 7432
rect 7607 7429 7619 7463
rect 7561 7423 7619 7429
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 8312 7460 8340 7500
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 11698 7528 11704 7540
rect 11563 7500 11704 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 11698 7488 11704 7500
rect 11756 7528 11762 7540
rect 12434 7528 12440 7540
rect 11756 7500 12440 7528
rect 11756 7488 11762 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 15286 7528 15292 7540
rect 13740 7500 14320 7528
rect 15247 7500 15292 7528
rect 8076 7432 8340 7460
rect 8076 7420 8082 7432
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 13740 7460 13768 7500
rect 9732 7432 13768 7460
rect 14292 7460 14320 7500
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 15930 7528 15936 7540
rect 15887 7500 15936 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 15930 7488 15936 7500
rect 15988 7528 15994 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15988 7500 16129 7528
rect 15988 7488 15994 7500
rect 16117 7497 16129 7500
rect 16163 7528 16175 7531
rect 16390 7528 16396 7540
rect 16163 7500 16396 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16390 7488 16396 7500
rect 16448 7528 16454 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16448 7500 16681 7528
rect 16448 7488 16454 7500
rect 16669 7497 16681 7500
rect 16715 7528 16727 7531
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16715 7500 17049 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 17678 7528 17684 7540
rect 17451 7500 17684 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 17052 7460 17080 7491
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 18012 7500 19073 7528
rect 18012 7488 18018 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 19061 7491 19119 7497
rect 21177 7531 21235 7537
rect 21177 7497 21189 7531
rect 21223 7528 21235 7531
rect 21358 7528 21364 7540
rect 21223 7500 21364 7528
rect 21223 7497 21235 7500
rect 21177 7491 21235 7497
rect 19518 7460 19524 7472
rect 14292 7432 16436 7460
rect 17052 7432 18828 7460
rect 9732 7420 9738 7432
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1636 7364 1869 7392
rect 1636 7352 1642 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 2314 7392 2320 7404
rect 2275 7364 2320 7392
rect 1857 7355 1915 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2464 7364 2789 7392
rect 2464 7352 2470 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3292 7364 4077 7392
rect 3292 7352 3298 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 4304 7364 5733 7392
rect 4304 7352 4310 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 8294 7392 8300 7404
rect 6420 7364 7880 7392
rect 8255 7364 8300 7392
rect 6420 7352 6426 7364
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 4798 7324 4804 7336
rect 3927 7296 4660 7324
rect 4759 7296 4804 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 1670 7216 1676 7268
rect 1728 7256 1734 7268
rect 1854 7256 1860 7268
rect 1728 7228 1860 7256
rect 1728 7216 1734 7228
rect 1854 7216 1860 7228
rect 1912 7216 1918 7268
rect 2958 7256 2964 7268
rect 2919 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 4632 7256 4660 7296
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 4982 7324 4988 7336
rect 4943 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 7006 7324 7012 7336
rect 6503 7296 7012 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7742 7324 7748 7336
rect 7703 7296 7748 7324
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7852 7324 7880 7364
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7392 11115 7395
rect 12066 7392 12072 7404
rect 11103 7364 12072 7392
rect 11103 7361 11115 7364
rect 11057 7355 11115 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12618 7392 12624 7404
rect 12676 7401 12682 7404
rect 12588 7364 12624 7392
rect 12618 7352 12624 7364
rect 12676 7355 12688 7401
rect 12676 7352 12682 7355
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12860 7364 12909 7392
rect 12860 7352 12866 7364
rect 12897 7361 12909 7364
rect 12943 7392 12955 7395
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 12943 7364 13185 7392
rect 12943 7361 12955 7364
rect 12897 7355 12955 7361
rect 13173 7361 13185 7364
rect 13219 7392 13231 7395
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 13219 7364 13553 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13541 7361 13553 7364
rect 13587 7392 13599 7395
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13587 7364 13921 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 14165 7395 14223 7401
rect 14165 7392 14177 7395
rect 13909 7355 13967 7361
rect 14016 7364 14177 7392
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 7852 7296 8585 7324
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 9398 7324 9404 7336
rect 9359 7296 9404 7324
rect 8573 7287 8631 7293
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7324 10011 7327
rect 10134 7324 10140 7336
rect 9999 7296 10140 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 14016 7324 14044 7364
rect 14165 7361 14177 7364
rect 14211 7361 14223 7395
rect 16408 7392 16436 7432
rect 17678 7392 17684 7404
rect 16408 7364 17684 7392
rect 14165 7355 14223 7361
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 18800 7401 18828 7432
rect 18892 7432 19524 7460
rect 18529 7395 18587 7401
rect 18529 7361 18541 7395
rect 18575 7392 18587 7395
rect 18785 7395 18843 7401
rect 18575 7364 18736 7392
rect 18575 7361 18587 7364
rect 18529 7355 18587 7361
rect 13188 7296 14044 7324
rect 18708 7324 18736 7364
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 18892 7324 18920 7432
rect 19518 7420 19524 7432
rect 19576 7460 19582 7472
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 19576 7432 20729 7460
rect 19576 7420 19582 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 20717 7423 20775 7429
rect 20174 7395 20232 7401
rect 20174 7392 20186 7395
rect 18708 7296 18920 7324
rect 19444 7364 20186 7392
rect 13188 7268 13216 7296
rect 5166 7256 5172 7268
rect 4632 7228 5172 7256
rect 5166 7216 5172 7228
rect 5224 7256 5230 7268
rect 5224 7228 10732 7256
rect 5224 7216 5230 7228
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7708 7160 8125 7188
rect 7708 7148 7714 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8113 7151 8171 7157
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 8260 7160 8953 7188
rect 8260 7148 8266 7160
rect 8941 7157 8953 7160
rect 8987 7157 8999 7191
rect 10226 7188 10232 7200
rect 10187 7160 10232 7188
rect 8941 7151 8999 7157
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10468 7160 10609 7188
rect 10468 7148 10474 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 10704 7188 10732 7228
rect 13170 7216 13176 7268
rect 13228 7216 13234 7268
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 19444 7256 19472 7364
rect 20174 7361 20186 7364
rect 20220 7361 20232 7395
rect 20174 7355 20232 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 21192 7392 21220 7491
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 20487 7364 21220 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 16264 7228 17908 7256
rect 16264 7216 16270 7228
rect 16758 7188 16764 7200
rect 10704 7160 16764 7188
rect 10597 7151 10655 7157
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 17880 7188 17908 7228
rect 18984 7228 19564 7256
rect 18984 7188 19012 7228
rect 19536 7200 19564 7228
rect 17880 7160 19012 7188
rect 19518 7148 19524 7200
rect 19576 7148 19582 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2682 6984 2688 6996
rect 2280 6956 2688 6984
rect 2280 6944 2286 6956
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 5040 6956 5181 6984
rect 5040 6944 5046 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 6822 6984 6828 6996
rect 5169 6947 5227 6953
rect 5552 6956 6828 6984
rect 4154 6916 4160 6928
rect 3896 6888 4160 6916
rect 2222 6848 2228 6860
rect 2183 6820 2228 6848
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 3896 6857 3924 6888
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 4890 6876 4896 6928
rect 4948 6916 4954 6928
rect 5552 6916 5580 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8352 6956 8953 6984
rect 8352 6944 8358 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 16206 6984 16212 6996
rect 8941 6947 8999 6953
rect 9048 6956 16212 6984
rect 4948 6888 5580 6916
rect 4948 6876 4954 6888
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 9048 6916 9076 6956
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 16390 6984 16396 6996
rect 16351 6956 16396 6984
rect 16390 6944 16396 6956
rect 16448 6984 16454 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 16448 6956 18429 6984
rect 16448 6944 16454 6956
rect 5684 6888 9076 6916
rect 9140 6888 9720 6916
rect 5684 6876 5690 6888
rect 3881 6851 3939 6857
rect 2832 6820 3556 6848
rect 2832 6808 2838 6820
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6780 1458 6792
rect 3418 6780 3424 6792
rect 1452 6752 3424 6780
rect 1452 6740 1458 6752
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 3528 6780 3556 6820
rect 3881 6817 3893 6851
rect 3927 6817 3939 6851
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 3881 6811 3939 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 5828 6857 5856 6888
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6817 5871 6851
rect 5813 6811 5871 6817
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 6880 6820 6925 6848
rect 7208 6820 7788 6848
rect 6880 6808 6886 6820
rect 6362 6780 6368 6792
rect 3528 6752 6368 6780
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 7208 6780 7236 6820
rect 7760 6789 7788 6820
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9140 6848 9168 6888
rect 8260 6820 9168 6848
rect 9585 6851 9643 6857
rect 8260 6808 8266 6820
rect 9585 6817 9597 6851
rect 9631 6817 9643 6851
rect 9692 6848 9720 6888
rect 13170 6876 13176 6928
rect 13228 6916 13234 6928
rect 13357 6919 13415 6925
rect 13357 6916 13369 6919
rect 13228 6888 13369 6916
rect 13228 6876 13234 6888
rect 13357 6885 13369 6888
rect 13403 6885 13415 6919
rect 13357 6879 13415 6885
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 9692 6820 10333 6848
rect 9585 6811 9643 6817
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 6687 6752 7236 6780
rect 7474 6776 7480 6788
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 7435 6748 7480 6776
rect 7474 6736 7480 6748
rect 7532 6736 7538 6788
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 9398 6780 9404 6792
rect 9355 6752 9404 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9600 6780 9628 6811
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11204 6820 11621 6848
rect 11204 6808 11210 6820
rect 11609 6817 11621 6820
rect 11655 6848 11667 6851
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11655 6820 11989 6848
rect 11655 6817 11667 6820
rect 11609 6811 11667 6817
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16408 6848 16436 6944
rect 18156 6860 18184 6956
rect 18417 6953 18429 6956
rect 18463 6984 18475 6987
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 18463 6956 18797 6984
rect 18463 6953 18475 6956
rect 18417 6947 18475 6953
rect 18785 6953 18797 6956
rect 18831 6984 18843 6987
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 18831 6956 19257 6984
rect 18831 6953 18843 6956
rect 18785 6947 18843 6953
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19613 6987 19671 6993
rect 19613 6984 19625 6987
rect 19576 6956 19625 6984
rect 19576 6944 19582 6956
rect 19613 6953 19625 6956
rect 19659 6953 19671 6987
rect 21358 6984 21364 6996
rect 19613 6947 19671 6953
rect 21008 6956 21364 6984
rect 21008 6860 21036 6956
rect 21358 6944 21364 6956
rect 21416 6944 21422 6996
rect 16080 6820 16436 6848
rect 16080 6808 16086 6820
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18196 6820 18289 6848
rect 18196 6808 18202 6820
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21048 6820 21141 6848
rect 21048 6808 21054 6820
rect 11698 6780 11704 6792
rect 9600 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12084 6752 15976 6780
rect 2409 6715 2467 6721
rect 2409 6681 2421 6715
rect 2455 6712 2467 6715
rect 3053 6715 3111 6721
rect 3053 6712 3065 6715
rect 2455 6684 3065 6712
rect 2455 6681 2467 6684
rect 2409 6675 2467 6681
rect 3053 6681 3065 6684
rect 3099 6681 3111 6715
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 3053 6675 3111 6681
rect 3528 6684 4169 6712
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2317 6647 2375 6653
rect 2317 6644 2329 6647
rect 1627 6616 2329 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2317 6613 2329 6616
rect 2363 6613 2375 6647
rect 2317 6607 2375 6613
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 3528 6644 3556 6684
rect 4157 6681 4169 6684
rect 4203 6681 4215 6715
rect 4801 6715 4859 6721
rect 4801 6712 4813 6715
rect 4157 6675 4215 6681
rect 4264 6684 4813 6712
rect 2823 6616 3556 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4264 6644 4292 6684
rect 4801 6681 4813 6684
rect 4847 6681 4859 6715
rect 4801 6675 4859 6681
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 5902 6712 5908 6724
rect 5583 6684 5908 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 10689 6715 10747 6721
rect 10689 6712 10701 6715
rect 7852 6684 10701 6712
rect 4522 6644 4528 6656
rect 4120 6616 4292 6644
rect 4483 6616 4528 6644
rect 4120 6604 4126 6616
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5224 6616 5641 6644
rect 5224 6604 5230 6616
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6273 6647 6331 6653
rect 6273 6644 6285 6647
rect 5776 6616 6285 6644
rect 5776 6604 5782 6616
rect 6273 6613 6285 6616
rect 6319 6613 6331 6647
rect 6273 6607 6331 6613
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 7282 6644 7288 6656
rect 6788 6616 6833 6644
rect 7243 6616 7288 6644
rect 6788 6604 6794 6616
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7852 6644 7880 6684
rect 10689 6681 10701 6684
rect 10735 6681 10747 6715
rect 10689 6675 10747 6681
rect 11333 6715 11391 6721
rect 11333 6681 11345 6715
rect 11379 6712 11391 6715
rect 12084 6712 12112 6752
rect 12233 6715 12291 6721
rect 12233 6712 12245 6715
rect 11379 6684 12112 6712
rect 12176 6684 12245 6712
rect 11379 6681 11391 6684
rect 11333 6675 11391 6681
rect 8294 6644 8300 6656
rect 7432 6616 7880 6644
rect 8255 6616 8300 6644
rect 7432 6604 7438 6616
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9088 6616 9413 6644
rect 9088 6604 9094 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9950 6644 9956 6656
rect 9911 6616 9956 6644
rect 9401 6607 9459 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 12176 6644 12204 6684
rect 12233 6681 12245 6684
rect 12279 6681 12291 6715
rect 12233 6675 12291 6681
rect 13725 6715 13783 6721
rect 13725 6681 13737 6715
rect 13771 6712 13783 6715
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 13771 6684 14381 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 14369 6681 14381 6684
rect 14415 6712 14427 6715
rect 15194 6712 15200 6724
rect 14415 6684 15200 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 15746 6672 15752 6724
rect 15804 6721 15810 6724
rect 15804 6712 15816 6721
rect 15948 6712 15976 6752
rect 17896 6715 17954 6721
rect 15804 6684 15849 6712
rect 15948 6684 17816 6712
rect 15804 6675 15816 6684
rect 15804 6672 15810 6675
rect 14642 6644 14648 6656
rect 11020 6616 12204 6644
rect 14603 6616 14648 6644
rect 11020 6604 11026 6616
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 16758 6644 16764 6656
rect 16719 6616 16764 6644
rect 16758 6604 16764 6616
rect 16816 6644 16822 6656
rect 17310 6644 17316 6656
rect 16816 6616 17316 6644
rect 16816 6604 16822 6616
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 17788 6644 17816 6684
rect 17896 6681 17908 6715
rect 17942 6712 17954 6715
rect 18046 6712 18052 6724
rect 17942 6684 18052 6712
rect 17942 6681 17954 6684
rect 17896 6675 17954 6681
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 19702 6672 19708 6724
rect 19760 6712 19766 6724
rect 20726 6715 20784 6721
rect 20726 6712 20738 6715
rect 19760 6684 20738 6712
rect 19760 6672 19766 6684
rect 20726 6681 20738 6684
rect 20772 6681 20784 6715
rect 20726 6675 20784 6681
rect 18322 6644 18328 6656
rect 17788 6616 18328 6644
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 19610 6644 19616 6656
rect 19024 6616 19616 6644
rect 19024 6604 19030 6616
rect 19610 6604 19616 6616
rect 19668 6604 19674 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 5534 6440 5540 6452
rect 4295 6412 5540 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5718 6440 5724 6452
rect 5675 6412 5724 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6454 6440 6460 6452
rect 6415 6412 6460 6440
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6730 6440 6736 6452
rect 6691 6412 6736 6440
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8168 6412 8585 6440
rect 8168 6400 8174 6412
rect 8573 6409 8585 6412
rect 8619 6440 8631 6443
rect 9030 6440 9036 6452
rect 8619 6412 8800 6440
rect 8991 6412 9036 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 8662 6372 8668 6384
rect 1412 6344 7236 6372
rect 8623 6344 8668 6372
rect 1412 6316 1440 6344
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 2832 6276 2877 6304
rect 2976 6276 3249 6304
rect 2832 6264 2838 6276
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2133 6239 2191 6245
rect 2133 6236 2145 6239
rect 1820 6208 2145 6236
rect 1820 6196 1826 6208
rect 2133 6205 2145 6208
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 2976 6236 3004 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 3326 6264 3332 6316
rect 3384 6304 3390 6316
rect 3605 6307 3663 6313
rect 3605 6304 3617 6307
rect 3384 6276 3617 6304
rect 3384 6264 3390 6276
rect 3605 6273 3617 6276
rect 3651 6273 3663 6307
rect 4062 6304 4068 6316
rect 3975 6276 4068 6304
rect 3605 6267 3663 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4580 6276 4813 6304
rect 4580 6264 4586 6276
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 7098 6304 7104 6316
rect 7059 6276 7104 6304
rect 4801 6267 4859 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7208 6304 7236 6344
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 8772 6372 8800 6412
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11204 6412 11529 6440
rect 11204 6400 11210 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 13170 6440 13176 6452
rect 11756 6412 13176 6440
rect 11756 6400 11762 6412
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6440 15531 6443
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 15519 6412 15853 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 15841 6409 15853 6412
rect 15887 6440 15899 6443
rect 16022 6440 16028 6452
rect 15887 6412 16028 6440
rect 15887 6409 15899 6412
rect 15841 6403 15899 6409
rect 9306 6372 9312 6384
rect 8772 6344 9312 6372
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 12802 6372 12808 6384
rect 10008 6344 12808 6372
rect 10008 6332 10014 6344
rect 12802 6332 12808 6344
rect 12860 6332 12866 6384
rect 13280 6344 15148 6372
rect 10226 6304 10232 6316
rect 7208 6276 10232 6304
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12158 6304 12164 6316
rect 11756 6276 12164 6304
rect 11756 6264 11762 6276
rect 12158 6264 12164 6276
rect 12216 6304 12222 6316
rect 12998 6307 13056 6313
rect 12998 6304 13010 6307
rect 12216 6276 13010 6304
rect 12216 6264 12222 6276
rect 12998 6273 13010 6276
rect 13044 6273 13056 6307
rect 12998 6267 13056 6273
rect 13170 6264 13176 6316
rect 13228 6264 13234 6316
rect 13280 6313 13308 6344
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6304 13323 6307
rect 13354 6304 13360 6316
rect 13311 6276 13360 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 14826 6264 14832 6316
rect 14884 6313 14890 6316
rect 15120 6313 15148 6344
rect 14884 6304 14896 6313
rect 15105 6307 15163 6313
rect 14884 6276 14929 6304
rect 14884 6267 14896 6276
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15194 6304 15200 6316
rect 15151 6276 15200 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 14884 6264 14890 6267
rect 15194 6264 15200 6276
rect 15252 6304 15258 6316
rect 15488 6304 15516 6403
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 16776 6412 18061 6440
rect 15252 6276 15516 6304
rect 16040 6304 16068 6400
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16040 6276 16681 6304
rect 15252 6264 15258 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 2924 6208 3004 6236
rect 2924 6196 2930 6208
rect 3050 6196 3056 6248
rect 3108 6236 3114 6248
rect 4080 6236 4108 6264
rect 3108 6208 4108 6236
rect 3108 6196 3114 6208
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5316 6208 5733 6236
rect 5316 6196 5322 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 2038 6168 2044 6180
rect 1627 6140 2044 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 2038 6128 2044 6140
rect 2096 6128 2102 6180
rect 4985 6171 5043 6177
rect 4985 6137 4997 6171
rect 5031 6168 5043 6171
rect 5626 6168 5632 6180
rect 5031 6140 5632 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 5828 6168 5856 6199
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 5960 6208 7205 6236
rect 5960 6196 5966 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7193 6199 7251 6205
rect 6454 6168 6460 6180
rect 5828 6140 6460 6168
rect 6454 6128 6460 6140
rect 6512 6128 6518 6180
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 7006 6168 7012 6180
rect 6604 6140 7012 6168
rect 6604 6128 6610 6140
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 7208 6168 7236 6199
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6205 8539 6239
rect 9306 6236 9312 6248
rect 9267 6208 9312 6236
rect 8481 6199 8539 6205
rect 7558 6168 7564 6180
rect 7208 6140 7564 6168
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 8496 6168 8524 6199
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 13188 6236 13216 6264
rect 13630 6236 13636 6248
rect 13188 6208 13636 6236
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 16776 6236 16804 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18064 6372 18092 6403
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 18196 6412 18337 6440
rect 18196 6400 18202 6412
rect 18325 6409 18337 6412
rect 18371 6440 18383 6443
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18371 6412 18705 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 18693 6409 18705 6412
rect 18739 6440 18751 6443
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18739 6412 19073 6440
rect 18739 6409 18751 6412
rect 18693 6403 18751 6409
rect 19061 6409 19073 6412
rect 19107 6440 19119 6443
rect 19107 6412 19196 6440
rect 19107 6409 19119 6412
rect 19061 6403 19119 6409
rect 18966 6372 18972 6384
rect 18064 6344 18972 6372
rect 18966 6332 18972 6344
rect 19024 6332 19030 6384
rect 16942 6313 16948 6316
rect 16936 6267 16948 6313
rect 17000 6304 17006 6316
rect 17000 6276 17036 6304
rect 16942 6264 16948 6267
rect 17000 6264 17006 6276
rect 17402 6264 17408 6316
rect 17460 6304 17466 6316
rect 19168 6304 19196 6412
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 20438 6440 20444 6452
rect 19300 6412 20444 6440
rect 19300 6400 19306 6412
rect 20438 6400 20444 6412
rect 20496 6440 20502 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 20496 6412 20821 6440
rect 20496 6400 20502 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 20809 6403 20867 6409
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 17460 6276 17724 6304
rect 19168 6276 19441 6304
rect 17460 6264 17466 6276
rect 16224 6208 16804 6236
rect 17696 6236 17724 6276
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 19685 6307 19743 6313
rect 19685 6304 19697 6307
rect 19429 6267 19487 6273
rect 19536 6276 19697 6304
rect 19536 6236 19564 6276
rect 19685 6273 19697 6276
rect 19731 6273 19743 6307
rect 19685 6267 19743 6273
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 21361 6307 21419 6313
rect 21361 6304 21373 6307
rect 21140 6276 21373 6304
rect 21140 6264 21146 6276
rect 21361 6273 21373 6276
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 17696 6208 19564 6236
rect 8496 6140 12112 6168
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 2593 6103 2651 6109
rect 2593 6100 2605 6103
rect 1728 6072 2605 6100
rect 1728 6060 1734 6072
rect 2593 6069 2605 6072
rect 2639 6069 2651 6103
rect 2593 6063 2651 6069
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6100 3111 6103
rect 3234 6100 3240 6112
rect 3099 6072 3240 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 4062 6100 4068 6112
rect 3835 6072 4068 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 4948 6072 5273 6100
rect 4948 6060 4954 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6730 6100 6736 6112
rect 5592 6072 6736 6100
rect 5592 6060 5598 6072
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 9490 6100 9496 6112
rect 8067 6072 9496 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10134 6100 10140 6112
rect 10095 6072 10140 6100
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10873 6103 10931 6109
rect 10873 6069 10885 6103
rect 10919 6100 10931 6103
rect 11790 6100 11796 6112
rect 10919 6072 11796 6100
rect 10919 6069 10931 6072
rect 10873 6063 10931 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12084 6100 12112 6140
rect 13722 6100 13728 6112
rect 11940 6072 11985 6100
rect 12084 6072 13728 6100
rect 11940 6060 11946 6072
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 16224 6100 16252 6208
rect 13872 6072 16252 6100
rect 16301 6103 16359 6109
rect 13872 6060 13878 6072
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 17586 6100 17592 6112
rect 16347 6072 17592 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 21174 6100 21180 6112
rect 21135 6072 21180 6100
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 2372 5868 3801 5896
rect 2372 5856 2378 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 5258 5896 5264 5908
rect 5219 5868 5264 5896
rect 3789 5859 3847 5865
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 6822 5896 6828 5908
rect 5368 5868 6828 5896
rect 2590 5788 2596 5840
rect 2648 5828 2654 5840
rect 3234 5828 3240 5840
rect 2648 5800 3240 5828
rect 2648 5788 2654 5800
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 1581 5763 1639 5769
rect 1581 5729 1593 5763
rect 1627 5760 1639 5763
rect 2501 5763 2559 5769
rect 2501 5760 2513 5763
rect 1627 5732 2513 5760
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 2501 5729 2513 5732
rect 2547 5760 2559 5763
rect 4522 5760 4528 5772
rect 2547 5732 4528 5760
rect 2547 5729 2559 5732
rect 2501 5723 2559 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4709 5763 4767 5769
rect 4709 5729 4721 5763
rect 4755 5760 4767 5763
rect 5368 5760 5396 5868
rect 6822 5856 6828 5868
rect 6880 5896 6886 5908
rect 8754 5896 8760 5908
rect 6880 5868 8760 5896
rect 6880 5856 6886 5868
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 8864 5868 9076 5896
rect 8294 5828 8300 5840
rect 6104 5800 8300 5828
rect 6104 5769 6132 5800
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 4755 5732 5396 5760
rect 6089 5763 6147 5769
rect 4755 5729 4767 5732
rect 4709 5723 4767 5729
rect 6089 5729 6101 5763
rect 6135 5729 6147 5763
rect 6089 5723 6147 5729
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 6512 5732 6929 5760
rect 6512 5720 6518 5732
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 8864 5760 8892 5868
rect 8941 5831 8999 5837
rect 8941 5797 8953 5831
rect 8987 5797 8999 5831
rect 9048 5828 9076 5868
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9858 5896 9864 5908
rect 9548 5868 9864 5896
rect 9548 5856 9554 5868
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10781 5899 10839 5905
rect 10781 5865 10793 5899
rect 10827 5896 10839 5899
rect 11146 5896 11152 5908
rect 10827 5868 11152 5896
rect 10827 5865 10839 5868
rect 10781 5859 10839 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 13354 5896 13360 5908
rect 11256 5868 13216 5896
rect 13315 5868 13360 5896
rect 11256 5828 11284 5868
rect 9048 5800 11284 5828
rect 13188 5828 13216 5868
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13630 5856 13636 5908
rect 13688 5896 13694 5908
rect 15841 5899 15899 5905
rect 13688 5868 15792 5896
rect 13688 5856 13694 5868
rect 14366 5828 14372 5840
rect 13188 5800 14372 5828
rect 8941 5791 8999 5797
rect 7515 5732 8892 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 3510 5692 3516 5704
rect 2823 5664 3516 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 4120 5664 7573 5692
rect 4120 5652 4126 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 7834 5692 7840 5704
rect 7699 5664 7840 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8956 5692 8984 5791
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 15764 5828 15792 5868
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16022 5896 16028 5908
rect 15887 5868 16028 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16022 5856 16028 5868
rect 16080 5896 16086 5908
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 16080 5868 16221 5896
rect 16080 5856 16086 5868
rect 16209 5865 16221 5868
rect 16255 5896 16267 5899
rect 16577 5899 16635 5905
rect 16577 5896 16589 5899
rect 16255 5868 16589 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 16577 5865 16589 5868
rect 16623 5865 16635 5899
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 16577 5859 16635 5865
rect 17052 5868 18429 5896
rect 17052 5828 17080 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 18417 5859 18475 5865
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 19702 5896 19708 5908
rect 19383 5868 19708 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 15764 5800 17080 5828
rect 18432 5828 18460 5859
rect 19702 5856 19708 5868
rect 19760 5856 19766 5908
rect 19794 5856 19800 5908
rect 19852 5856 19858 5908
rect 19812 5828 19840 5856
rect 18432 5800 19840 5828
rect 20990 5788 20996 5840
rect 21048 5788 21054 5840
rect 9030 5720 9036 5772
rect 9088 5760 9094 5772
rect 9585 5763 9643 5769
rect 9088 5732 9536 5760
rect 9088 5720 9094 5732
rect 9306 5692 9312 5704
rect 8527 5664 8984 5692
rect 9267 5664 9312 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 1670 5624 1676 5636
rect 1631 5596 1676 5624
rect 1670 5584 1676 5596
rect 1728 5584 1734 5636
rect 3234 5584 3240 5636
rect 3292 5624 3298 5636
rect 6181 5627 6239 5633
rect 6181 5624 6193 5627
rect 3292 5596 6193 5624
rect 3292 5584 3298 5596
rect 6181 5593 6193 5596
rect 6227 5593 6239 5627
rect 7926 5624 7932 5636
rect 6181 5587 6239 5593
rect 6656 5596 7932 5624
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5556 2191 5559
rect 2406 5556 2412 5568
rect 2179 5528 2412 5556
rect 2179 5525 2191 5528
rect 2133 5519 2191 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2685 5559 2743 5565
rect 2685 5525 2697 5559
rect 2731 5556 2743 5559
rect 2958 5556 2964 5568
rect 2731 5528 2964 5556
rect 2731 5525 2743 5528
rect 2685 5519 2743 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 3602 5556 3608 5568
rect 3191 5528 3608 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4798 5556 4804 5568
rect 4759 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 4893 5559 4951 5565
rect 4893 5525 4905 5559
rect 4939 5556 4951 5559
rect 5166 5556 5172 5568
rect 4939 5528 5172 5556
rect 4939 5525 4951 5528
rect 4893 5519 4951 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 6656 5565 6684 5596
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8036 5596 9413 5624
rect 8036 5565 8064 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9508 5624 9536 5732
rect 9585 5729 9597 5763
rect 9631 5729 9643 5763
rect 9585 5723 9643 5729
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 13354 5760 13360 5772
rect 12851 5732 13360 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 9600 5692 9628 5723
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 14458 5760 14464 5772
rect 13648 5732 14464 5760
rect 13648 5692 13676 5732
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 16022 5760 16028 5772
rect 15519 5732 16028 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 16022 5720 16028 5732
rect 16080 5760 16086 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16080 5732 17049 5760
rect 16080 5720 16086 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5760 20775 5763
rect 21008 5760 21036 5788
rect 20763 5732 21036 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 9600 5664 13676 5692
rect 13722 5652 13728 5704
rect 13780 5692 13786 5704
rect 17293 5695 17351 5701
rect 17293 5692 17305 5695
rect 13780 5664 17305 5692
rect 13780 5652 13786 5664
rect 17293 5661 17305 5664
rect 17339 5661 17351 5695
rect 17293 5655 17351 5661
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 18693 5695 18751 5701
rect 18693 5692 18705 5695
rect 17644 5664 18705 5692
rect 17644 5652 17650 5664
rect 18693 5661 18705 5664
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 12560 5627 12618 5633
rect 9508 5596 12434 5624
rect 9401 5587 9459 5593
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 5776 5528 6285 5556
rect 5776 5516 5782 5528
rect 6273 5525 6285 5528
rect 6319 5525 6331 5559
rect 6273 5519 6331 5525
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5525 6699 5559
rect 6641 5519 6699 5525
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5525 8079 5559
rect 8294 5556 8300 5568
rect 8255 5528 8300 5556
rect 8021 5519 8079 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 9950 5556 9956 5568
rect 9911 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 11020 5528 11437 5556
rect 11020 5516 11026 5528
rect 11425 5525 11437 5528
rect 11471 5525 11483 5559
rect 12406 5556 12434 5596
rect 12560 5593 12572 5627
rect 12606 5624 12618 5627
rect 14274 5624 14280 5636
rect 12606 5596 14280 5624
rect 12606 5593 12618 5596
rect 12560 5587 12618 5593
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 15228 5627 15286 5633
rect 15228 5593 15240 5627
rect 15274 5624 15286 5627
rect 15562 5624 15568 5636
rect 15274 5596 15568 5624
rect 15274 5593 15286 5596
rect 15228 5587 15286 5593
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 15746 5584 15752 5636
rect 15804 5624 15810 5636
rect 17954 5624 17960 5636
rect 15804 5596 17960 5624
rect 15804 5584 15810 5596
rect 17954 5584 17960 5596
rect 18012 5584 18018 5636
rect 18708 5624 18736 5655
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 19484 5664 21005 5692
rect 19484 5652 19490 5664
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 20070 5624 20076 5636
rect 18708 5596 20076 5624
rect 20070 5584 20076 5596
rect 20128 5584 20134 5636
rect 20438 5584 20444 5636
rect 20496 5633 20502 5636
rect 20496 5624 20508 5633
rect 20496 5596 20541 5624
rect 20496 5587 20508 5596
rect 20496 5584 20502 5587
rect 13814 5556 13820 5568
rect 12406 5528 13820 5556
rect 11425 5519 11483 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 18230 5556 18236 5568
rect 14424 5528 18236 5556
rect 14424 5516 14430 5528
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 18877 5559 18935 5565
rect 18877 5525 18889 5559
rect 18923 5556 18935 5559
rect 19242 5556 19248 5568
rect 18923 5528 19248 5556
rect 18923 5525 18935 5528
rect 18877 5519 18935 5525
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 20772 5528 21189 5556
rect 20772 5516 20778 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 21177 5519 21235 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2590 5352 2596 5364
rect 2551 5324 2596 5352
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 2958 5352 2964 5364
rect 2919 5324 2964 5352
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3237 5355 3295 5361
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 3510 5352 3516 5364
rect 3283 5324 3516 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 4062 5352 4068 5364
rect 3743 5324 4068 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4798 5352 4804 5364
rect 4755 5324 4804 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5258 5352 5264 5364
rect 5215 5324 5264 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5258 5312 5264 5324
rect 5316 5352 5322 5364
rect 5902 5352 5908 5364
rect 5316 5324 5908 5352
rect 5316 5312 5322 5324
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 6546 5352 6552 5364
rect 6144 5324 6552 5352
rect 6144 5312 6150 5324
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 8110 5352 8116 5364
rect 6779 5324 8116 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 3605 5287 3663 5293
rect 3605 5284 3617 5287
rect 3476 5256 3617 5284
rect 3476 5244 3482 5256
rect 3605 5253 3617 5256
rect 3651 5284 3663 5287
rect 6748 5284 6776 5315
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9950 5352 9956 5364
rect 9171 5324 9956 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 11882 5352 11888 5364
rect 10152 5324 11888 5352
rect 3651 5256 4752 5284
rect 3651 5253 3663 5256
rect 3605 5247 3663 5253
rect 4724 5228 4752 5256
rect 5552 5256 6776 5284
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 2498 5216 2504 5228
rect 2459 5188 2504 5216
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 4246 5216 4252 5228
rect 3068 5188 3832 5216
rect 4207 5188 4252 5216
rect 1412 5080 1440 5176
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 3068 5148 3096 5188
rect 3804 5160 3832 5188
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4706 5176 4712 5228
rect 4764 5176 4770 5228
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 4856 5188 5089 5216
rect 4856 5176 4862 5188
rect 5077 5185 5089 5188
rect 5123 5216 5135 5219
rect 5552 5216 5580 5256
rect 7926 5244 7932 5296
rect 7984 5284 7990 5296
rect 9217 5287 9275 5293
rect 9217 5284 9229 5287
rect 7984 5256 9229 5284
rect 7984 5244 7990 5256
rect 9217 5253 9229 5256
rect 9263 5253 9275 5287
rect 9217 5247 9275 5253
rect 5123 5188 5580 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5684 5188 5733 5216
rect 5684 5176 5690 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7561 5219 7619 5225
rect 6871 5188 7052 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 2455 5120 3096 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3602 5148 3608 5160
rect 3200 5120 3608 5148
rect 3200 5108 3206 5120
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 3786 5148 3792 5160
rect 3747 5120 3792 5148
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 5350 5148 5356 5160
rect 5311 5120 5356 5148
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6840 5148 6868 5179
rect 5960 5120 6868 5148
rect 6917 5151 6975 5157
rect 5960 5108 5966 5120
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 7024 5148 7052 5188
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8478 5216 8484 5228
rect 7607 5188 8484 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 10042 5216 10048 5228
rect 8588 5188 10048 5216
rect 8588 5148 8616 5188
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 7024 5120 8616 5148
rect 6917 5111 6975 5117
rect 5258 5080 5264 5092
rect 1412 5052 5264 5080
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 6730 5040 6736 5092
rect 6788 5080 6794 5092
rect 6932 5080 6960 5111
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9122 5148 9128 5160
rect 8720 5120 9128 5148
rect 8720 5108 8726 5120
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 10152 5148 10180 5324
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 13265 5355 13323 5361
rect 12575 5324 13216 5352
rect 10904 5287 10962 5293
rect 10904 5253 10916 5287
rect 10950 5284 10962 5287
rect 12575 5284 12603 5324
rect 10950 5256 12603 5284
rect 13188 5284 13216 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5352 13418 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13412 5324 13553 5352
rect 13412 5312 13418 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 16209 5355 16267 5361
rect 16209 5352 16221 5355
rect 16080 5324 16221 5352
rect 16080 5312 16086 5324
rect 16209 5321 16221 5324
rect 16255 5321 16267 5355
rect 19426 5352 19432 5364
rect 19387 5324 19432 5352
rect 16209 5315 16267 5321
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 13188 5256 15893 5284
rect 10950 5253 10962 5256
rect 10904 5247 10962 5253
rect 11146 5216 11152 5228
rect 11107 5188 11152 5216
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 12618 5176 12624 5228
rect 12676 5225 12682 5228
rect 12676 5216 12688 5225
rect 12897 5219 12955 5225
rect 12676 5188 12721 5216
rect 12676 5179 12688 5188
rect 12897 5185 12909 5219
rect 12943 5216 12955 5219
rect 13354 5216 13360 5228
rect 12943 5188 13360 5216
rect 12943 5185 12955 5188
rect 12897 5179 12955 5185
rect 12676 5176 12682 5179
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 15666 5219 15724 5225
rect 15666 5216 15678 5219
rect 14148 5188 15678 5216
rect 14148 5176 14154 5188
rect 15666 5185 15678 5188
rect 15712 5185 15724 5219
rect 15666 5179 15724 5185
rect 11698 5148 11704 5160
rect 9447 5120 10180 5148
rect 11532 5120 11704 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 11532 5089 11560 5120
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 15865 5148 15893 5256
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16040 5216 16068 5312
rect 16936 5287 16994 5293
rect 16936 5253 16948 5287
rect 16982 5284 16994 5287
rect 17126 5284 17132 5296
rect 16982 5256 17132 5284
rect 16982 5253 16994 5256
rect 16936 5247 16994 5253
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 21174 5284 21180 5296
rect 17236 5256 21180 5284
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 15979 5188 16681 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 17236 5216 17264 5256
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 16669 5179 16727 5185
rect 16776 5188 17264 5216
rect 16776 5148 16804 5188
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18693 5219 18751 5225
rect 18693 5216 18705 5219
rect 18564 5188 18705 5216
rect 18564 5176 18570 5188
rect 18693 5185 18705 5188
rect 18739 5185 18751 5219
rect 19242 5216 19248 5228
rect 19203 5188 19248 5216
rect 18693 5179 18751 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 20806 5216 20812 5228
rect 20864 5225 20870 5228
rect 20776 5188 20812 5216
rect 20806 5176 20812 5188
rect 20864 5179 20876 5225
rect 20864 5176 20870 5179
rect 20990 5176 20996 5228
rect 21048 5216 21054 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 21048 5188 21097 5216
rect 21048 5176 21054 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 15865 5120 16804 5148
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 18104 5120 19748 5148
rect 18104 5108 18110 5120
rect 6788 5052 6960 5080
rect 8481 5083 8539 5089
rect 6788 5040 6794 5052
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 11517 5083 11575 5089
rect 8527 5052 9444 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 9416 5024 9444 5052
rect 11517 5049 11529 5083
rect 11563 5049 11575 5083
rect 18325 5083 18383 5089
rect 18325 5080 18337 5083
rect 11517 5043 11575 5049
rect 17604 5052 18337 5080
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 5012 1918 5024
rect 3970 5012 3976 5024
rect 1912 4984 3976 5012
rect 1912 4972 1918 4984
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 4982 5012 4988 5024
rect 4479 4984 4988 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 4982 4972 4988 4984
rect 5040 5012 5046 5024
rect 5626 5012 5632 5024
rect 5040 4984 5632 5012
rect 5040 4972 5046 4984
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 5902 5012 5908 5024
rect 5863 4984 5908 5012
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 7064 4984 7389 5012
rect 7064 4972 7070 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 7377 4975 7435 4981
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 8628 4984 8769 5012
rect 8628 4972 8634 4984
rect 8757 4981 8769 4984
rect 8803 4981 8815 5015
rect 8757 4975 8815 4981
rect 9398 4972 9404 5024
rect 9456 4972 9462 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 5012 9827 5015
rect 9950 5012 9956 5024
rect 9815 4984 9956 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 11756 4984 13921 5012
rect 11756 4972 11762 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 14550 5012 14556 5024
rect 14511 4984 14556 5012
rect 13909 4975 13967 4981
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 17604 5012 17632 5052
rect 18325 5049 18337 5052
rect 18371 5080 18383 5083
rect 18506 5080 18512 5092
rect 18371 5052 18512 5080
rect 18371 5049 18383 5052
rect 18325 5043 18383 5049
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 19720 5089 19748 5120
rect 19705 5083 19763 5089
rect 19705 5049 19717 5083
rect 19751 5049 19763 5083
rect 19705 5043 19763 5049
rect 15804 4984 17632 5012
rect 18049 5015 18107 5021
rect 15804 4972 15810 4984
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18138 5012 18144 5024
rect 18095 4984 18144 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18656 4984 18889 5012
rect 18656 4972 18662 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 18877 4975 18935 4981
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 4525 4811 4583 4817
rect 2608 4780 3280 4808
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 2130 4672 2136 4684
rect 1995 4644 2136 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4672 2283 4675
rect 2608 4672 2636 4780
rect 3142 4700 3148 4752
rect 3200 4700 3206 4752
rect 3252 4740 3280 4780
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4614 4808 4620 4820
rect 4571 4780 4620 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 12621 4811 12679 4817
rect 6880 4780 9628 4808
rect 6880 4768 6886 4780
rect 3252 4712 8524 4740
rect 2271 4644 2636 4672
rect 2685 4675 2743 4681
rect 2271 4641 2283 4644
rect 2225 4635 2283 4641
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 2958 4672 2964 4684
rect 2731 4644 2964 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 2240 4604 2268 4635
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 1912 4576 2268 4604
rect 1912 4564 1918 4576
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2464 4576 2881 4604
rect 2464 4564 2470 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 3160 4536 3188 4700
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6362 4672 6368 4684
rect 5767 4644 6368 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4604 4123 4607
rect 4430 4604 4436 4616
rect 4111 4576 4436 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5258 4604 5264 4616
rect 5215 4576 5264 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 2823 4508 3188 4536
rect 4724 4536 4752 4567
rect 5258 4564 5264 4576
rect 5316 4604 5322 4616
rect 5534 4604 5540 4616
rect 5316 4576 5540 4604
rect 5316 4564 5322 4576
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5644 4604 5672 4635
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 8386 4672 8392 4684
rect 7331 4644 8392 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 6730 4604 6736 4616
rect 5644 4576 6736 4604
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7650 4604 7656 4616
rect 7611 4576 7656 4604
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8294 4604 8300 4616
rect 8255 4576 8300 4604
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8496 4604 8524 4712
rect 9600 4681 9628 4780
rect 12621 4777 12633 4811
rect 12667 4808 12679 4811
rect 12894 4808 12900 4820
rect 12667 4780 12900 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 13354 4808 13360 4820
rect 13035 4780 13360 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13354 4768 13360 4780
rect 13412 4808 13418 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13412 4780 13645 4808
rect 13412 4768 13418 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 14274 4768 14280 4820
rect 14332 4808 14338 4820
rect 14332 4780 17632 4808
rect 14332 4768 14338 4780
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 14737 4743 14795 4749
rect 14737 4740 14749 4743
rect 12584 4712 14749 4740
rect 12584 4700 12590 4712
rect 14737 4709 14749 4712
rect 14783 4709 14795 4743
rect 14737 4703 14795 4709
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 17497 4743 17555 4749
rect 17497 4740 17509 4743
rect 16356 4712 17509 4740
rect 16356 4700 16362 4712
rect 17497 4709 17509 4712
rect 17543 4709 17555 4743
rect 17497 4703 17555 4709
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 10962 4672 10968 4684
rect 9815 4644 10968 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 11204 4644 11253 4672
rect 11204 4632 11210 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 16942 4672 16948 4684
rect 11241 4635 11299 4641
rect 16316 4644 16948 4672
rect 10318 4604 10324 4616
rect 8496 4576 10324 4604
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 11256 4604 11284 4635
rect 11256 4576 12434 4604
rect 12406 4548 12434 4576
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 14461 4607 14519 4613
rect 12860 4576 14412 4604
rect 12860 4564 12866 4576
rect 5350 4536 5356 4548
rect 4724 4508 5356 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 5350 4496 5356 4508
rect 5408 4536 5414 4548
rect 6086 4536 6092 4548
rect 5408 4508 6092 4536
rect 5408 4496 5414 4508
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 7101 4539 7159 4545
rect 7101 4536 7113 4539
rect 6196 4508 7113 4536
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 5074 4468 5080 4480
rect 5031 4440 5080 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 6196 4477 6224 4508
rect 7101 4505 7113 4508
rect 7147 4505 7159 4539
rect 7101 4499 7159 4505
rect 8496 4508 10916 4536
rect 6181 4471 6239 4477
rect 5868 4440 5913 4468
rect 5868 4428 5874 4440
rect 6181 4437 6193 4471
rect 6227 4437 6239 4471
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6181 4431 6239 4437
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7009 4471 7067 4477
rect 7009 4437 7021 4471
rect 7055 4468 7067 4471
rect 7374 4468 7380 4480
rect 7055 4440 7380 4468
rect 7055 4437 7067 4440
rect 7009 4431 7067 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7834 4468 7840 4480
rect 7795 4440 7840 4468
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 8496 4477 8524 4508
rect 8481 4471 8539 4477
rect 8481 4437 8493 4471
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 8904 4440 9137 4468
rect 8904 4428 8910 4440
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 9490 4468 9496 4480
rect 9451 4440 9496 4468
rect 9125 4431 9183 4437
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 9732 4440 10149 4468
rect 9732 4428 9738 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10888 4468 10916 4508
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 11238 4536 11244 4548
rect 11112 4508 11244 4536
rect 11112 4496 11118 4508
rect 11238 4496 11244 4508
rect 11296 4536 11302 4548
rect 11486 4539 11544 4545
rect 11486 4536 11498 4539
rect 11296 4508 11498 4536
rect 11296 4496 11302 4508
rect 11486 4505 11498 4508
rect 11532 4505 11544 4539
rect 11486 4499 11544 4505
rect 12342 4496 12348 4548
rect 12400 4536 12434 4548
rect 13354 4536 13360 4548
rect 12400 4508 13360 4536
rect 12400 4496 12406 4508
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 14384 4536 14412 4576
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 14507 4576 15976 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 15746 4536 15752 4548
rect 14384 4508 15752 4536
rect 15746 4496 15752 4508
rect 15804 4536 15810 4548
rect 15850 4539 15908 4545
rect 15850 4536 15862 4539
rect 15804 4508 15862 4536
rect 15804 4496 15810 4508
rect 15850 4505 15862 4508
rect 15896 4505 15908 4539
rect 15948 4536 15976 4576
rect 16022 4564 16028 4616
rect 16080 4604 16086 4616
rect 16117 4607 16175 4613
rect 16117 4604 16129 4607
rect 16080 4576 16129 4604
rect 16080 4564 16086 4576
rect 16117 4573 16129 4576
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 16316 4536 16344 4644
rect 16942 4632 16948 4644
rect 17000 4632 17006 4684
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 17604 4604 17632 4780
rect 18230 4768 18236 4820
rect 18288 4808 18294 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 18288 4780 19257 4808
rect 18288 4768 18294 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 19245 4771 19303 4777
rect 20625 4675 20683 4681
rect 20625 4641 20637 4675
rect 20671 4672 20683 4675
rect 20990 4672 20996 4684
rect 20671 4644 20996 4672
rect 20671 4641 20683 4644
rect 20625 4635 20683 4641
rect 18877 4607 18935 4613
rect 17604 4576 18736 4604
rect 16393 4567 16451 4573
rect 15948 4508 16344 4536
rect 15850 4499 15908 4505
rect 12434 4468 12440 4480
rect 10888 4440 12440 4468
rect 10137 4431 10195 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 13538 4428 13544 4480
rect 13596 4468 13602 4480
rect 14277 4471 14335 4477
rect 14277 4468 14289 4471
rect 13596 4440 14289 4468
rect 13596 4428 13602 4440
rect 14277 4437 14289 4440
rect 14323 4437 14335 4471
rect 14277 4431 14335 4437
rect 14366 4428 14372 4480
rect 14424 4468 14430 4480
rect 16408 4468 16436 4567
rect 18414 4536 18420 4548
rect 16592 4508 18420 4536
rect 16592 4477 16620 4508
rect 18414 4496 18420 4508
rect 18472 4496 18478 4548
rect 18610 4539 18668 4545
rect 18610 4536 18622 4539
rect 18524 4508 18622 4536
rect 14424 4440 16436 4468
rect 16577 4471 16635 4477
rect 14424 4428 14430 4440
rect 16577 4437 16589 4471
rect 16623 4437 16635 4471
rect 17034 4468 17040 4480
rect 16995 4440 17040 4468
rect 16577 4431 16635 4437
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18524 4468 18552 4508
rect 18610 4505 18622 4508
rect 18656 4505 18668 4539
rect 18610 4499 18668 4505
rect 17920 4440 18552 4468
rect 18708 4468 18736 4576
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 20640 4604 20668 4635
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 18923 4576 20668 4604
rect 20901 4607 20959 4613
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19720 4548 19748 4576
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21450 4604 21456 4616
rect 20947 4576 21456 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21450 4564 21456 4576
rect 21508 4564 21514 4616
rect 19702 4496 19708 4548
rect 19760 4496 19766 4548
rect 20358 4539 20416 4545
rect 20358 4536 20370 4539
rect 19812 4508 20370 4536
rect 19812 4468 19840 4508
rect 20358 4505 20370 4508
rect 20404 4505 20416 4539
rect 20358 4499 20416 4505
rect 21082 4468 21088 4480
rect 18708 4440 19840 4468
rect 21043 4440 21088 4468
rect 17920 4428 17926 4440
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 3513 4267 3571 4273
rect 3513 4264 3525 4267
rect 3476 4236 3525 4264
rect 3476 4224 3482 4236
rect 3513 4233 3525 4236
rect 3559 4233 3571 4267
rect 3513 4227 3571 4233
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 7558 4264 7564 4276
rect 4304 4236 7564 4264
rect 4304 4224 4310 4236
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 8941 4267 8999 4273
rect 8941 4233 8953 4267
rect 8987 4233 8999 4267
rect 8941 4227 8999 4233
rect 11701 4267 11759 4273
rect 11701 4233 11713 4267
rect 11747 4264 11759 4267
rect 12158 4264 12164 4276
rect 11747 4236 12164 4264
rect 11747 4233 11759 4236
rect 11701 4227 11759 4233
rect 4338 4196 4344 4208
rect 3804 4168 4344 4196
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1820 4100 1961 4128
rect 1820 4088 1826 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 1949 4091 2007 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 3234 4128 3240 4140
rect 2731 4100 3240 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3804 4137 3832 4168
rect 4338 4156 4344 4168
rect 4396 4196 4402 4208
rect 4982 4196 4988 4208
rect 4396 4168 4988 4196
rect 4396 4156 4402 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 5537 4199 5595 4205
rect 5537 4165 5549 4199
rect 5583 4196 5595 4199
rect 5626 4196 5632 4208
rect 5583 4168 5632 4196
rect 5583 4165 5595 4168
rect 5537 4159 5595 4165
rect 5626 4156 5632 4168
rect 5684 4196 5690 4208
rect 6178 4196 6184 4208
rect 5684 4168 6184 4196
rect 5684 4156 5690 4168
rect 6178 4156 6184 4168
rect 6236 4156 6242 4208
rect 6914 4156 6920 4208
rect 6972 4156 6978 4208
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 3344 4060 3372 4091
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 4154 4128 4160 4140
rect 3936 4100 4160 4128
rect 3936 4088 3942 4100
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4709 4131 4767 4137
rect 4304 4100 4349 4128
rect 4304 4088 4310 4100
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 5074 4128 5080 4140
rect 4755 4100 5080 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 6270 4128 6276 4140
rect 5644 4100 6276 4128
rect 4062 4060 4068 4072
rect 3344 4032 4068 4060
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 5644 4069 5672 4100
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6457 4131 6515 4137
rect 6457 4097 6469 4131
rect 6503 4128 6515 4131
rect 6932 4128 6960 4156
rect 6503 4100 6960 4128
rect 6503 4097 6515 4100
rect 6457 4091 6515 4097
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7248 4100 7389 4128
rect 7248 4088 7254 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7650 4128 7656 4140
rect 7524 4100 7656 4128
rect 7524 4088 7530 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8956 4128 8984 4227
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12342 4264 12348 4276
rect 12303 4236 12348 4264
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 15102 4264 15108 4276
rect 12492 4236 15108 4264
rect 12492 4224 12498 4236
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 16850 4264 16856 4276
rect 15580 4236 16856 4264
rect 9309 4199 9367 4205
rect 9309 4165 9321 4199
rect 9355 4196 9367 4199
rect 9674 4196 9680 4208
rect 9355 4168 9680 4196
rect 9355 4165 9367 4168
rect 9309 4159 9367 4165
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 10796 4168 11652 4196
rect 8711 4100 8984 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 5902 4060 5908 4072
rect 5859 4032 5908 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6914 4060 6920 4072
rect 6875 4032 6920 4060
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 8036 4060 8064 4091
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9766 4128 9772 4140
rect 9180 4100 9772 4128
rect 9180 4088 9186 4100
rect 9766 4088 9772 4100
rect 9824 4128 9830 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 9824 4100 10149 4128
rect 9824 4088 9830 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10796 4128 10824 4168
rect 10744 4100 10824 4128
rect 10744 4088 10750 4100
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 10928 4100 11161 4128
rect 10928 4088 10934 4100
rect 11149 4097 11161 4100
rect 11195 4097 11207 4131
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11149 4091 11207 4097
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11624 4128 11652 4168
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 13412 4168 13860 4196
rect 13412 4156 13418 4168
rect 11624 4100 13032 4128
rect 7024 4032 8064 4060
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 3602 3992 3608 4004
rect 3292 3964 3608 3992
rect 3292 3952 3298 3964
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 3970 3992 3976 4004
rect 3931 3964 3976 3992
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4430 3992 4436 4004
rect 4391 3964 4436 3992
rect 4430 3952 4436 3964
rect 4488 3952 4494 4004
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 4893 3995 4951 4001
rect 4893 3992 4905 3995
rect 4856 3964 4905 3992
rect 4856 3952 4862 3964
rect 4893 3961 4905 3964
rect 4939 3961 4951 3995
rect 5166 3992 5172 4004
rect 5127 3964 5172 3992
rect 4893 3955 4951 3961
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 7024 3992 7052 4032
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 9401 4063 9459 4069
rect 9401 4060 9413 4063
rect 8904 4032 9413 4060
rect 8904 4020 8910 4032
rect 9401 4029 9413 4032
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4029 9551 4063
rect 12894 4060 12900 4072
rect 9493 4023 9551 4029
rect 10060 4032 12900 4060
rect 5592 3964 7052 3992
rect 7561 3995 7619 4001
rect 5592 3952 5598 3964
rect 7561 3961 7573 3995
rect 7607 3992 7619 3995
rect 7607 3964 8892 3992
rect 7607 3961 7619 3964
rect 7561 3955 7619 3961
rect 2869 3927 2927 3933
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 3418 3924 3424 3936
rect 2915 3896 3424 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 8018 3924 8024 3936
rect 6687 3896 8024 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8478 3924 8484 3936
rect 8439 3896 8484 3924
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8864 3924 8892 3964
rect 9306 3952 9312 4004
rect 9364 3992 9370 4004
rect 9508 3992 9536 4023
rect 9950 3992 9956 4004
rect 9364 3964 9536 3992
rect 9911 3964 9956 3992
rect 9364 3952 9370 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10060 3924 10088 4032
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 10689 3995 10747 4001
rect 10689 3961 10701 3995
rect 10735 3992 10747 3995
rect 11054 3992 11060 4004
rect 10735 3964 11060 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 11054 3952 11060 3964
rect 11112 3992 11118 4004
rect 11514 3992 11520 4004
rect 11112 3964 11520 3992
rect 11112 3952 11118 3964
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3992 12679 3995
rect 12802 3992 12808 4004
rect 12667 3964 12808 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 8864 3896 10088 3924
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 10965 3927 11023 3933
rect 10965 3924 10977 3927
rect 10560 3896 10977 3924
rect 10560 3884 10566 3896
rect 10965 3893 10977 3896
rect 11011 3893 11023 3927
rect 10965 3887 11023 3893
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11882 3924 11888 3936
rect 11388 3896 11888 3924
rect 11388 3884 11394 3896
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 13004 3924 13032 4100
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13734 4131 13792 4137
rect 13734 4128 13746 4131
rect 13320 4100 13746 4128
rect 13320 4088 13326 4100
rect 13734 4097 13746 4100
rect 13780 4097 13792 4131
rect 13832 4128 13860 4168
rect 14458 4156 14464 4208
rect 14516 4196 14522 4208
rect 15580 4196 15608 4236
rect 16850 4224 16856 4236
rect 16908 4264 16914 4276
rect 17862 4264 17868 4276
rect 16908 4236 17868 4264
rect 16908 4224 16914 4236
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 16022 4196 16028 4208
rect 14516 4168 15608 4196
rect 15672 4168 16028 4196
rect 14516 4156 14522 4168
rect 15672 4137 15700 4168
rect 16022 4156 16028 4168
rect 16080 4156 16086 4208
rect 20990 4156 20996 4208
rect 21048 4196 21054 4208
rect 21048 4168 21404 4196
rect 21048 4156 21054 4168
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13832 4100 14013 4128
rect 13734 4091 13792 4097
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 15401 4131 15459 4137
rect 15401 4097 15413 4131
rect 15447 4128 15459 4131
rect 15657 4131 15715 4137
rect 15447 4100 15608 4128
rect 15447 4097 15459 4100
rect 15401 4091 15459 4097
rect 15580 4060 15608 4100
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15930 4128 15936 4140
rect 15891 4100 15936 4128
rect 15657 4091 15715 4097
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 16040 4128 16068 4156
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16040 4100 16681 4128
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16936 4131 16994 4137
rect 16936 4097 16948 4131
rect 16982 4128 16994 4131
rect 17218 4128 17224 4140
rect 16982 4100 17224 4128
rect 16982 4097 16994 4100
rect 16936 4091 16994 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 19426 4088 19432 4140
rect 19484 4137 19490 4140
rect 19484 4128 19496 4137
rect 19702 4128 19708 4140
rect 19484 4100 19529 4128
rect 19663 4100 19708 4128
rect 19484 4091 19496 4100
rect 19484 4088 19490 4091
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 21105 4131 21163 4137
rect 21105 4097 21117 4131
rect 21151 4128 21163 4131
rect 21266 4128 21272 4140
rect 21151 4100 21272 4128
rect 21151 4097 21163 4100
rect 21105 4091 21163 4097
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 21376 4137 21404 4168
rect 21361 4131 21419 4137
rect 21361 4097 21373 4131
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 15580 4032 16528 4060
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 13004 3896 14289 3924
rect 14277 3893 14289 3896
rect 14323 3893 14335 3927
rect 14277 3887 14335 3893
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16390 3924 16396 3936
rect 16163 3896 16396 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 16500 3924 16528 4032
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18325 3995 18383 4001
rect 18325 3992 18337 3995
rect 18012 3964 18337 3992
rect 18012 3952 18018 3964
rect 18325 3961 18337 3964
rect 18371 3961 18383 3995
rect 18325 3955 18383 3961
rect 17310 3924 17316 3936
rect 16500 3896 17316 3924
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17828 3896 18061 3924
rect 17828 3884 17834 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 18564 3896 19993 3924
rect 18564 3884 18570 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 19981 3887 20039 3893
rect 1104 3834 21896 3856
rect 14 3748 20 3800
rect 72 3788 78 3800
rect 934 3788 940 3800
rect 72 3760 940 3788
rect 72 3748 78 3760
rect 934 3748 940 3760
rect 992 3748 998 3800
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 4706 3720 4712 3732
rect 4663 3692 4712 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5534 3720 5540 3732
rect 5495 3692 5540 3720
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5810 3720 5816 3732
rect 5771 3692 5816 3720
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 6822 3720 6828 3732
rect 6328 3692 6828 3720
rect 6328 3680 6334 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 8352 3692 8401 3720
rect 8352 3680 8358 3692
rect 8389 3689 8401 3692
rect 8435 3689 8447 3723
rect 8389 3683 8447 3689
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 15930 3720 15936 3732
rect 8904 3692 15936 3720
rect 8904 3680 8910 3692
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 16945 3723 17003 3729
rect 16945 3720 16957 3723
rect 16908 3692 16957 3720
rect 16908 3680 16914 3692
rect 16945 3689 16957 3692
rect 16991 3689 17003 3723
rect 16945 3683 17003 3689
rect 17236 3692 18368 3720
rect 5077 3655 5135 3661
rect 5077 3621 5089 3655
rect 5123 3652 5135 3655
rect 5123 3624 8708 3652
rect 5123 3621 5135 3624
rect 5077 3615 5135 3621
rect 8680 3596 8708 3624
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 9309 3655 9367 3661
rect 9309 3652 9321 3655
rect 8996 3624 9321 3652
rect 8996 3612 9002 3624
rect 9309 3621 9321 3624
rect 9355 3621 9367 3655
rect 9309 3615 9367 3621
rect 9585 3655 9643 3661
rect 9585 3621 9597 3655
rect 9631 3652 9643 3655
rect 9766 3652 9772 3664
rect 9631 3624 9772 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 11241 3655 11299 3661
rect 11241 3621 11253 3655
rect 11287 3652 11299 3655
rect 11330 3652 11336 3664
rect 11287 3624 11336 3652
rect 11287 3621 11299 3624
rect 11241 3615 11299 3621
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 14093 3655 14151 3661
rect 14093 3621 14105 3655
rect 14139 3652 14151 3655
rect 14274 3652 14280 3664
rect 14139 3624 14280 3652
rect 14139 3621 14151 3624
rect 14093 3615 14151 3621
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 15562 3612 15568 3664
rect 15620 3652 15626 3664
rect 16577 3655 16635 3661
rect 15620 3624 16160 3652
rect 15620 3612 15626 3624
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2958 3544 2964 3596
rect 3016 3584 3022 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 3016 3556 3341 3584
rect 3016 3544 3022 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 6086 3584 6092 3596
rect 3329 3547 3387 3553
rect 4448 3556 6092 3584
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 992 3488 2237 3516
rect 992 3476 998 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3234 3516 3240 3528
rect 3099 3488 3240 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 4448 3525 4476 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6270 3584 6276 3596
rect 6231 3556 6276 3584
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6546 3584 6552 3596
rect 6503 3556 6552 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6546 3544 6552 3556
rect 6604 3584 6610 3596
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 6604 3556 7665 3584
rect 6604 3544 6610 3556
rect 7653 3553 7665 3556
rect 7699 3553 7711 3587
rect 7653 3547 7711 3553
rect 7834 3544 7840 3596
rect 7892 3584 7898 3596
rect 8110 3584 8116 3596
rect 7892 3556 8116 3584
rect 7892 3544 7898 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8662 3544 8668 3596
rect 8720 3544 8726 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9674 3584 9680 3596
rect 9456 3556 9680 3584
rect 9456 3544 9462 3556
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11146 3584 11152 3596
rect 11011 3556 11152 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 16022 3584 16028 3596
rect 15519 3556 16028 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 16132 3584 16160 3624
rect 16577 3621 16589 3655
rect 16623 3652 16635 3655
rect 17126 3652 17132 3664
rect 16623 3624 17132 3652
rect 16623 3621 16635 3624
rect 16577 3615 16635 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 17236 3584 17264 3692
rect 18340 3652 18368 3692
rect 18966 3680 18972 3732
rect 19024 3720 19030 3732
rect 21082 3720 21088 3732
rect 19024 3692 21088 3720
rect 19024 3680 19030 3692
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 19245 3655 19303 3661
rect 19245 3652 19257 3655
rect 18340 3624 19257 3652
rect 19245 3621 19257 3624
rect 19291 3621 19303 3655
rect 19245 3615 19303 3621
rect 16132 3556 17264 3584
rect 18325 3587 18383 3593
rect 18325 3553 18337 3587
rect 18371 3584 18383 3587
rect 18506 3584 18512 3596
rect 18371 3556 18512 3584
rect 18371 3553 18383 3556
rect 18325 3547 18383 3553
rect 18506 3544 18512 3556
rect 18564 3584 18570 3596
rect 19610 3584 19616 3596
rect 18564 3556 19616 3584
rect 18564 3544 18570 3556
rect 19610 3544 19616 3556
rect 19668 3544 19674 3596
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3476 3488 3985 3516
rect 3476 3476 3482 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4890 3516 4896 3528
rect 4851 3488 4896 3516
rect 4433 3479 4491 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 6638 3516 6644 3528
rect 5399 3488 6644 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7466 3516 7472 3528
rect 7427 3488 7472 3516
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 8570 3516 8576 3528
rect 7616 3488 7661 3516
rect 8531 3488 8576 3516
rect 7616 3476 7622 3488
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 10226 3516 10232 3528
rect 9600 3504 10232 3516
rect 9125 3479 9183 3485
rect 5442 3448 5448 3460
rect 4172 3420 5448 3448
rect 4172 3389 4200 3420
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 6086 3408 6092 3460
rect 6144 3448 6150 3460
rect 6546 3448 6552 3460
rect 6144 3420 6552 3448
rect 6144 3408 6150 3420
rect 6546 3408 6552 3420
rect 6604 3408 6610 3460
rect 9582 3452 9588 3504
rect 9640 3488 10232 3504
rect 9640 3452 9646 3488
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10686 3476 10692 3528
rect 10744 3525 10750 3528
rect 10744 3516 10756 3525
rect 11164 3516 11192 3544
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 10744 3488 10789 3516
rect 11164 3488 12633 3516
rect 10744 3479 10756 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3485 12955 3519
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 12897 3479 12955 3485
rect 10744 3476 10750 3479
rect 10778 3408 10784 3460
rect 10836 3448 10842 3460
rect 12354 3451 12412 3457
rect 12354 3448 12366 3451
rect 10836 3420 12366 3448
rect 10836 3408 10842 3420
rect 12354 3417 12366 3420
rect 12400 3448 12412 3451
rect 12526 3448 12532 3460
rect 12400 3420 12532 3448
rect 12400 3417 12412 3420
rect 12354 3411 12412 3417
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3349 4215 3383
rect 4157 3343 4215 3349
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 5902 3380 5908 3392
rect 5316 3352 5908 3380
rect 5316 3340 5322 3352
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 6178 3380 6184 3392
rect 6139 3352 6184 3380
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 7098 3380 7104 3392
rect 7059 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 9490 3340 9496 3392
rect 9548 3380 9554 3392
rect 12912 3380 12940 3479
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 15206 3519 15264 3525
rect 15206 3516 15218 3519
rect 14700 3488 15218 3516
rect 14700 3476 14706 3488
rect 15206 3485 15218 3488
rect 15252 3485 15264 3519
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 15206 3479 15264 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18472 3488 18613 3516
rect 18472 3476 18478 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 19628 3516 19656 3544
rect 20530 3516 20536 3528
rect 19628 3488 20536 3516
rect 18601 3479 18659 3485
rect 20530 3476 20536 3488
rect 20588 3516 20594 3528
rect 20625 3519 20683 3525
rect 20625 3516 20637 3519
rect 20588 3488 20637 3516
rect 20588 3476 20594 3488
rect 20625 3485 20637 3488
rect 20671 3485 20683 3519
rect 20625 3479 20683 3485
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3516 20959 3519
rect 20990 3516 20996 3528
rect 20947 3488 20996 3516
rect 20947 3485 20959 3488
rect 20901 3479 20959 3485
rect 20990 3476 20996 3488
rect 21048 3476 21054 3528
rect 15010 3448 15016 3460
rect 13096 3420 15016 3448
rect 13096 3389 13124 3420
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 18138 3457 18144 3460
rect 18080 3451 18144 3457
rect 18080 3417 18092 3451
rect 18126 3417 18144 3451
rect 18080 3411 18144 3417
rect 18138 3408 18144 3411
rect 18196 3408 18202 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 18288 3420 19380 3448
rect 18288 3408 18294 3420
rect 9548 3352 12940 3380
rect 13081 3383 13139 3389
rect 9548 3340 9554 3352
rect 13081 3349 13093 3383
rect 13127 3349 13139 3383
rect 13081 3343 13139 3349
rect 13725 3383 13783 3389
rect 13725 3349 13737 3383
rect 13771 3380 13783 3383
rect 13814 3380 13820 3392
rect 13771 3352 13820 3380
rect 13771 3349 13783 3352
rect 13725 3343 13783 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 16025 3383 16083 3389
rect 16025 3349 16037 3383
rect 16071 3380 16083 3383
rect 16390 3380 16396 3392
rect 16071 3352 16396 3380
rect 16071 3349 16083 3352
rect 16025 3343 16083 3349
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 17552 3352 18797 3380
rect 17552 3340 17558 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 19352 3380 19380 3420
rect 19794 3408 19800 3460
rect 19852 3448 19858 3460
rect 20358 3451 20416 3457
rect 20358 3448 20370 3451
rect 19852 3420 20370 3448
rect 19852 3408 19858 3420
rect 20358 3417 20370 3420
rect 20404 3417 20416 3451
rect 20358 3411 20416 3417
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 19352 3352 21097 3380
rect 18785 3343 18843 3349
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 5074 3176 5080 3188
rect 5035 3148 5080 3176
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5534 3176 5540 3188
rect 5495 3148 5540 3176
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6972 3148 7021 3176
rect 6972 3136 6978 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7374 3176 7380 3188
rect 7335 3148 7380 3176
rect 7009 3139 7067 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8110 3176 8116 3188
rect 8071 3148 8116 3176
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8573 3179 8631 3185
rect 8573 3145 8585 3179
rect 8619 3176 8631 3179
rect 8846 3176 8852 3188
rect 8619 3148 8852 3176
rect 8619 3145 8631 3148
rect 8573 3139 8631 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9033 3179 9091 3185
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9306 3176 9312 3188
rect 9079 3148 9312 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9490 3176 9496 3188
rect 9451 3148 9496 3176
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 12400 3148 13369 3176
rect 12400 3136 12406 3148
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 13357 3139 13415 3145
rect 15013 3179 15071 3185
rect 15013 3145 15025 3179
rect 15059 3145 15071 3179
rect 15013 3139 15071 3145
rect 16669 3179 16727 3185
rect 16669 3145 16681 3179
rect 16715 3176 16727 3179
rect 16850 3176 16856 3188
rect 16715 3148 16856 3176
rect 16715 3145 16727 3148
rect 16669 3139 16727 3145
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 7282 3108 7288 3120
rect 2648 3080 2774 3108
rect 2648 3068 2654 3080
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1544 3012 1961 3040
rect 1544 3000 1550 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 2746 3040 2774 3080
rect 5828 3080 7288 3108
rect 3234 3040 3240 3052
rect 2746 3012 3240 3040
rect 1949 3003 2007 3009
rect 3234 3000 3240 3012
rect 3292 3040 3298 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3292 3012 3617 3040
rect 3292 3000 3298 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 5828 3049 5856 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 8938 3068 8944 3120
rect 8996 3108 9002 3120
rect 8996 3080 12434 3108
rect 8996 3068 9002 3080
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3752 3012 3893 3040
rect 3752 3000 3758 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5813 3043 5871 3049
rect 5399 3012 5764 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2774 2972 2780 2984
rect 2271 2944 2780 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 3142 2972 3148 2984
rect 3099 2944 3148 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3418 2972 3424 2984
rect 3375 2944 3424 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 4908 2972 4936 3003
rect 5736 2972 5764 3012
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 7098 3040 7104 3052
rect 6963 3012 7104 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 8386 3040 8392 3052
rect 8347 3012 8392 3040
rect 7929 3003 7987 3009
rect 6730 2972 6736 2984
rect 4908 2944 5672 2972
rect 5736 2944 6132 2972
rect 6691 2944 6736 2972
rect 5644 2836 5672 2944
rect 5994 2904 6000 2916
rect 5955 2876 6000 2904
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 6104 2904 6132 2944
rect 6730 2932 6736 2944
rect 6788 2972 6794 2984
rect 7834 2972 7840 2984
rect 6788 2944 7840 2972
rect 6788 2932 6794 2944
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 7944 2972 7972 3003
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 9214 3040 9220 3052
rect 8849 3027 8907 3033
rect 8849 2993 8861 3027
rect 8895 3024 8907 3027
rect 8956 3024 9220 3040
rect 8895 3012 9220 3024
rect 8895 2996 8984 3012
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9674 3040 9680 3052
rect 9355 3012 9680 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9674 3000 9680 3012
rect 9732 3040 9738 3052
rect 10502 3040 10508 3052
rect 9732 3012 10508 3040
rect 9732 3000 9738 3012
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 10882 3043 10940 3049
rect 10882 3040 10894 3043
rect 10652 3012 10894 3040
rect 10652 3000 10658 3012
rect 10882 3009 10894 3012
rect 10928 3009 10940 3043
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 10882 3003 10940 3009
rect 11146 3000 11152 3012
rect 11204 3040 11210 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11204 3012 11529 3040
rect 11204 3000 11210 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11773 3043 11831 3049
rect 11773 3040 11785 3043
rect 11517 3003 11575 3009
rect 11624 3012 11785 3040
rect 8895 2993 8907 2996
rect 8849 2987 8907 2993
rect 8662 2972 8668 2984
rect 7944 2944 8668 2972
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 9232 2972 9260 3000
rect 9766 2972 9772 2984
rect 9232 2944 9772 2972
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 11624 2972 11652 3012
rect 11773 3009 11785 3012
rect 11819 3009 11831 3043
rect 12406 3040 12434 3080
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 15028 3108 15056 3139
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17034 3176 17040 3188
rect 16995 3148 17040 3176
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 21266 3176 21272 3188
rect 17920 3148 21272 3176
rect 17920 3136 17926 3148
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 12952 3080 14872 3108
rect 15028 3080 17724 3108
rect 12952 3068 12958 3080
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 12406 3012 13185 3040
rect 11773 3003 11831 3009
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13722 3040 13728 3052
rect 13683 3012 13728 3040
rect 13173 3003 13231 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14844 3049 14872 3080
rect 14277 3043 14335 3049
rect 14277 3009 14289 3043
rect 14323 3009 14335 3043
rect 14277 3003 14335 3009
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 14829 3003 14887 3009
rect 11532 2944 11652 2972
rect 7558 2904 7564 2916
rect 6104 2876 7564 2904
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8018 2864 8024 2916
rect 8076 2904 8082 2916
rect 9214 2904 9220 2916
rect 8076 2876 9220 2904
rect 8076 2864 8082 2876
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 7190 2836 7196 2848
rect 5644 2808 7196 2836
rect 7190 2796 7196 2808
rect 7248 2836 7254 2848
rect 7650 2836 7656 2848
rect 7248 2808 7656 2836
rect 7248 2796 7254 2808
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 7800 2808 9781 2836
rect 7800 2796 7806 2808
rect 9769 2805 9781 2808
rect 9815 2836 9827 2839
rect 11532 2836 11560 2944
rect 13354 2932 13360 2984
rect 13412 2972 13418 2984
rect 14292 2972 14320 3003
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15930 3040 15936 3052
rect 15891 3012 15936 3040
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 17696 3049 17724 3080
rect 18322 3068 18328 3120
rect 18380 3108 18386 3120
rect 18380 3080 20208 3108
rect 18380 3068 18386 3080
rect 17681 3043 17739 3049
rect 16960 3012 17632 3040
rect 13412 2944 14320 2972
rect 13412 2932 13418 2944
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 16960 2972 16988 3012
rect 14424 2944 16988 2972
rect 14424 2932 14430 2944
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 17092 2944 17141 2972
rect 17092 2932 17098 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2941 17371 2975
rect 17604 2972 17632 3012
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 17681 3003 17739 3009
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 20180 3049 20208 3080
rect 18765 3043 18823 3049
rect 18765 3040 18777 3043
rect 18616 3012 18777 3040
rect 17770 2972 17776 2984
rect 17604 2944 17776 2972
rect 17313 2935 17371 2941
rect 12897 2907 12955 2913
rect 12897 2873 12909 2907
rect 12943 2904 12955 2907
rect 13262 2904 13268 2916
rect 12943 2876 13268 2904
rect 12943 2873 12955 2876
rect 12897 2867 12955 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 17328 2904 17356 2935
rect 17770 2932 17776 2944
rect 17828 2972 17834 2984
rect 18616 2972 18644 3012
rect 18765 3009 18777 3012
rect 18811 3009 18823 3043
rect 18765 3003 18823 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3040 20223 3043
rect 20806 3040 20812 3052
rect 20211 3012 20812 3040
rect 20211 3009 20223 3012
rect 20165 3003 20223 3009
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 20530 2972 20536 2984
rect 17828 2944 18644 2972
rect 20491 2944 20536 2972
rect 17828 2932 17834 2944
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 17328 2876 18552 2904
rect 9815 2808 11560 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 13446 2796 13452 2848
rect 13504 2836 13510 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 13504 2808 13921 2836
rect 13504 2796 13510 2808
rect 13909 2805 13921 2808
rect 13955 2805 13967 2839
rect 13909 2799 13967 2805
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 14332 2808 14473 2836
rect 14332 2796 14338 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 15565 2839 15623 2845
rect 15565 2836 15577 2839
rect 15344 2808 15577 2836
rect 15344 2796 15350 2808
rect 15565 2805 15577 2808
rect 15611 2805 15623 2839
rect 15565 2799 15623 2805
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 16117 2839 16175 2845
rect 16117 2836 16129 2839
rect 15712 2808 16129 2836
rect 15712 2796 15718 2808
rect 16117 2805 16129 2808
rect 16163 2805 16175 2839
rect 16117 2799 16175 2805
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 17865 2839 17923 2845
rect 17865 2836 17877 2839
rect 17000 2808 17877 2836
rect 17000 2796 17006 2808
rect 17865 2805 17877 2808
rect 17911 2805 17923 2839
rect 18524 2836 18552 2876
rect 19518 2836 19524 2848
rect 18524 2808 19524 2836
rect 17865 2799 17923 2805
rect 19518 2796 19524 2808
rect 19576 2836 19582 2848
rect 19889 2839 19947 2845
rect 19889 2836 19901 2839
rect 19576 2808 19901 2836
rect 19576 2796 19582 2808
rect 19889 2805 19901 2808
rect 19935 2805 19947 2839
rect 19889 2799 19947 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 11146 2632 11152 2644
rect 9079 2604 11152 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 11146 2592 11152 2604
rect 11204 2632 11210 2644
rect 11204 2604 12940 2632
rect 11204 2592 11210 2604
rect 2498 2564 2504 2576
rect 1964 2536 2504 2564
rect 1964 2505 1992 2536
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 4798 2524 4804 2576
rect 4856 2524 4862 2576
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 6638 2564 6644 2576
rect 6043 2536 6644 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 6638 2524 6644 2536
rect 6696 2524 6702 2576
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 9214 2564 9220 2576
rect 8619 2536 9220 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 9858 2564 9864 2576
rect 9416 2536 9864 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 2314 2496 2320 2508
rect 2271 2468 2320 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2038 2388 2044 2440
rect 2096 2428 2102 2440
rect 2240 2428 2268 2459
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 2464 2468 3341 2496
rect 2464 2456 2470 2468
rect 3329 2465 3341 2468
rect 3375 2496 3387 2499
rect 3970 2496 3976 2508
rect 3375 2468 3976 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 3970 2456 3976 2468
rect 4028 2456 4034 2508
rect 4816 2496 4844 2524
rect 7098 2496 7104 2508
rect 4264 2468 4844 2496
rect 4908 2468 7104 2496
rect 2096 2400 2268 2428
rect 3053 2431 3111 2437
rect 2096 2388 2102 2400
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 4264 2428 4292 2468
rect 3099 2400 4292 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4617 2431 4675 2437
rect 4396 2400 4441 2428
rect 4396 2388 4402 2400
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 4798 2428 4804 2440
rect 4663 2400 4804 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 4908 2437 4936 2468
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 8478 2496 8484 2508
rect 7484 2468 8484 2496
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 5534 2428 5540 2440
rect 5399 2400 5540 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6822 2428 6828 2440
rect 6595 2400 6828 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 7006 2428 7012 2440
rect 6967 2400 7012 2428
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7484 2437 7512 2468
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7926 2428 7932 2440
rect 7887 2400 7932 2428
rect 7469 2391 7527 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 9416 2428 9444 2536
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 11238 2524 11244 2576
rect 11296 2564 11302 2576
rect 11517 2567 11575 2573
rect 11517 2564 11529 2567
rect 11296 2536 11529 2564
rect 11296 2524 11302 2536
rect 11517 2533 11529 2536
rect 11563 2533 11575 2567
rect 11517 2527 11575 2533
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2496 9551 2499
rect 11790 2496 11796 2508
rect 9539 2468 9996 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 8435 2400 9444 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9732 2400 9777 2428
rect 9732 2388 9738 2400
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 4246 2360 4252 2372
rect 4120 2332 4252 2360
rect 4120 2320 4126 2332
rect 4246 2320 4252 2332
rect 4304 2360 4310 2372
rect 9600 2360 9628 2388
rect 4304 2332 9628 2360
rect 9968 2360 9996 2468
rect 10520 2468 11796 2496
rect 10520 2437 10548 2468
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12912 2505 12940 2604
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 19334 2632 19340 2644
rect 16632 2604 19340 2632
rect 16632 2592 16638 2604
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 19702 2632 19708 2644
rect 19444 2604 19708 2632
rect 13078 2524 13084 2576
rect 13136 2564 13142 2576
rect 14277 2567 14335 2573
rect 14277 2564 14289 2567
rect 13136 2536 14289 2564
rect 13136 2524 13142 2536
rect 14277 2533 14289 2536
rect 14323 2533 14335 2567
rect 14277 2527 14335 2533
rect 14550 2524 14556 2576
rect 14608 2564 14614 2576
rect 15381 2567 15439 2573
rect 15381 2564 15393 2567
rect 14608 2536 15393 2564
rect 14608 2524 14614 2536
rect 15381 2533 15393 2536
rect 15427 2533 15439 2567
rect 15381 2527 15439 2533
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 17405 2567 17463 2573
rect 17405 2564 17417 2567
rect 16448 2536 17417 2564
rect 16448 2524 16454 2536
rect 17405 2533 17417 2536
rect 17451 2533 17463 2567
rect 17405 2527 17463 2533
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 13872 2468 14688 2496
rect 13872 2456 13878 2468
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 11698 2428 11704 2440
rect 11195 2400 11704 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 12641 2431 12699 2437
rect 12641 2397 12653 2431
rect 12687 2428 12699 2431
rect 12802 2428 12808 2440
rect 12687 2400 12808 2428
rect 12687 2397 12699 2400
rect 12641 2391 12699 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 13170 2428 13176 2440
rect 13131 2400 13176 2428
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14660 2437 14688 2468
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 18049 2499 18107 2505
rect 15160 2468 15792 2496
rect 15160 2456 15166 2468
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 14645 2391 14703 2397
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15764 2437 15792 2468
rect 18049 2465 18061 2499
rect 18095 2496 18107 2499
rect 19444 2496 19472 2604
rect 19702 2592 19708 2604
rect 19760 2632 19766 2644
rect 20162 2632 20168 2644
rect 19760 2604 20168 2632
rect 19760 2592 19766 2604
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 21266 2632 21272 2644
rect 21227 2604 21272 2632
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 18095 2468 19472 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 15838 2388 15844 2440
rect 15896 2428 15902 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 15896 2400 16681 2428
rect 15896 2388 15902 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 17221 2391 17279 2397
rect 9968 2332 13492 2360
rect 4304 2320 4310 2332
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 5077 2295 5135 2301
rect 5077 2292 5089 2295
rect 1360 2264 5089 2292
rect 1360 2252 1366 2264
rect 5077 2261 5089 2264
rect 5123 2261 5135 2295
rect 5077 2255 5135 2261
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2292 5595 2295
rect 5902 2292 5908 2304
rect 5583 2264 5908 2292
rect 5583 2261 5595 2264
rect 5537 2255 5595 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 6730 2292 6736 2304
rect 6691 2264 6736 2292
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 7193 2295 7251 2301
rect 7193 2261 7205 2295
rect 7239 2292 7251 2295
rect 7466 2292 7472 2304
rect 7239 2264 7472 2292
rect 7239 2261 7251 2264
rect 7193 2255 7251 2261
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 7650 2292 7656 2304
rect 7611 2264 7656 2292
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 9398 2292 9404 2304
rect 7984 2264 9404 2292
rect 7984 2252 7990 2264
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 9585 2295 9643 2301
rect 9585 2261 9597 2295
rect 9631 2292 9643 2295
rect 9674 2292 9680 2304
rect 9631 2264 9680 2292
rect 9631 2261 9643 2264
rect 9585 2255 9643 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10686 2292 10692 2304
rect 10647 2264 10692 2292
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 10962 2292 10968 2304
rect 10923 2264 10968 2292
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 12860 2264 13369 2292
rect 12860 2252 12866 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13464 2292 13492 2332
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 13872 2332 14872 2360
rect 13872 2320 13878 2332
rect 14366 2292 14372 2304
rect 13464 2264 14372 2292
rect 13357 2255 13415 2261
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 14844 2301 14872 2332
rect 15010 2320 15016 2372
rect 15068 2360 15074 2372
rect 17236 2360 17264 2391
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 19518 2428 19524 2440
rect 19475 2400 19524 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2428 21143 2431
rect 21450 2428 21456 2440
rect 21131 2400 21456 2428
rect 21131 2397 21143 2400
rect 21085 2391 21143 2397
rect 21450 2388 21456 2400
rect 21508 2388 21514 2440
rect 15068 2332 17264 2360
rect 15068 2320 15074 2332
rect 18138 2320 18144 2372
rect 18196 2360 18202 2372
rect 19674 2363 19732 2369
rect 19674 2360 19686 2363
rect 18196 2332 19686 2360
rect 18196 2320 18202 2332
rect 19674 2329 19686 2332
rect 19720 2329 19732 2363
rect 19674 2323 19732 2329
rect 14829 2295 14887 2301
rect 14829 2261 14841 2295
rect 14875 2261 14887 2295
rect 14829 2255 14887 2261
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 15933 2295 15991 2301
rect 15933 2292 15945 2295
rect 14976 2264 15945 2292
rect 14976 2252 14982 2264
rect 15933 2261 15945 2264
rect 15979 2261 15991 2295
rect 15933 2255 15991 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16080 2264 16865 2292
rect 16080 2252 16086 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20772 2264 20821 2292
rect 20772 2252 20778 2264
rect 20809 2261 20821 2264
rect 20855 2292 20867 2295
rect 20898 2292 20904 2304
rect 20855 2264 20904 2292
rect 20855 2261 20867 2264
rect 20809 2255 20867 2261
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 5534 2048 5540 2100
rect 5592 2088 5598 2100
rect 8294 2088 8300 2100
rect 5592 2060 8300 2088
rect 5592 2048 5598 2060
rect 8294 2048 8300 2060
rect 8352 2048 8358 2100
rect 13170 2088 13176 2100
rect 9600 2060 13176 2088
rect 5442 1980 5448 2032
rect 5500 2020 5506 2032
rect 9600 2020 9628 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 5500 1992 9628 2020
rect 5500 1980 5506 1992
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 17034 2020 17040 2032
rect 10100 1992 17040 2020
rect 10100 1980 10106 1992
rect 17034 1980 17040 1992
rect 17092 1980 17098 2032
rect 7466 1912 7472 1964
rect 7524 1952 7530 1964
rect 15838 1952 15844 1964
rect 7524 1924 15844 1952
rect 7524 1912 7530 1924
rect 15838 1912 15844 1924
rect 15896 1912 15902 1964
rect 20714 1952 20720 1964
rect 16546 1924 20720 1952
rect 4062 1844 4068 1896
rect 4120 1884 4126 1896
rect 4798 1884 4804 1896
rect 4120 1856 4804 1884
rect 4120 1844 4126 1856
rect 4798 1844 4804 1856
rect 4856 1884 4862 1896
rect 10410 1884 10416 1896
rect 4856 1856 10416 1884
rect 4856 1844 4862 1856
rect 10410 1844 10416 1856
rect 10468 1844 10474 1896
rect 10686 1844 10692 1896
rect 10744 1884 10750 1896
rect 12434 1884 12440 1896
rect 10744 1856 12440 1884
rect 10744 1844 10750 1856
rect 12434 1844 12440 1856
rect 12492 1844 12498 1896
rect 5810 1776 5816 1828
rect 5868 1816 5874 1828
rect 8662 1816 8668 1828
rect 5868 1788 8668 1816
rect 5868 1776 5874 1788
rect 8662 1776 8668 1788
rect 8720 1776 8726 1828
rect 14090 1816 14096 1828
rect 11808 1788 14096 1816
rect 7834 1708 7840 1760
rect 7892 1748 7898 1760
rect 7892 1720 8064 1748
rect 7892 1708 7898 1720
rect 7098 1640 7104 1692
rect 7156 1680 7162 1692
rect 7926 1680 7932 1692
rect 7156 1652 7932 1680
rect 7156 1640 7162 1652
rect 7926 1640 7932 1652
rect 7984 1640 7990 1692
rect 8036 1680 8064 1720
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 11808 1748 11836 1788
rect 14090 1776 14096 1788
rect 14148 1776 14154 1828
rect 8260 1720 11836 1748
rect 8260 1708 8266 1720
rect 12066 1708 12072 1760
rect 12124 1748 12130 1760
rect 15378 1748 15384 1760
rect 12124 1720 15384 1748
rect 12124 1708 12130 1720
rect 15378 1708 15384 1720
rect 15436 1708 15442 1760
rect 16546 1748 16574 1924
rect 20714 1912 20720 1924
rect 20772 1912 20778 1964
rect 15488 1720 16574 1748
rect 15488 1680 15516 1720
rect 18322 1680 18328 1692
rect 8036 1652 15516 1680
rect 16546 1652 18328 1680
rect 11606 1572 11612 1624
rect 11664 1612 11670 1624
rect 11790 1612 11796 1624
rect 11664 1584 11796 1612
rect 11664 1572 11670 1584
rect 11790 1572 11796 1584
rect 11848 1572 11854 1624
rect 16546 1612 16574 1652
rect 18322 1640 18328 1652
rect 18380 1640 18386 1692
rect 12406 1584 16574 1612
rect 5718 1504 5724 1556
rect 5776 1544 5782 1556
rect 6454 1544 6460 1556
rect 5776 1516 6460 1544
rect 5776 1504 5782 1516
rect 6454 1504 6460 1516
rect 6512 1504 6518 1556
rect 7650 1436 7656 1488
rect 7708 1476 7714 1488
rect 12066 1476 12072 1488
rect 7708 1448 12072 1476
rect 7708 1436 7714 1448
rect 12066 1436 12072 1448
rect 12124 1436 12130 1488
rect 9674 1368 9680 1420
rect 9732 1408 9738 1420
rect 9950 1408 9956 1420
rect 9732 1380 9956 1408
rect 9732 1368 9738 1380
rect 9950 1368 9956 1380
rect 10008 1408 10014 1420
rect 12406 1408 12434 1584
rect 10008 1380 12434 1408
rect 10008 1368 10014 1380
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 2780 20544 2832 20596
rect 4436 20408 4488 20460
rect 1860 20340 1912 20392
rect 2964 20340 3016 20392
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 2872 20000 2924 20052
rect 4436 20043 4488 20052
rect 4436 20009 4445 20043
rect 4445 20009 4479 20043
rect 4479 20009 4488 20043
rect 4436 20000 4488 20009
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 10416 19796 10468 19848
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 2228 19456 2280 19508
rect 5724 19456 5776 19508
rect 1952 19320 2004 19372
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 7288 19320 7340 19372
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 2044 19227 2096 19236
rect 2044 19193 2053 19227
rect 2053 19193 2087 19227
rect 2087 19193 2096 19227
rect 2044 19184 2096 19193
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1676 18912 1728 18964
rect 3884 18708 3936 18760
rect 5908 18708 5960 18760
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 2228 18368 2280 18420
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 7472 18232 7524 18284
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1676 17824 1728 17876
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 5908 17824 5960 17876
rect 1952 17756 2004 17808
rect 1952 17620 2004 17672
rect 2596 17620 2648 17672
rect 3608 17552 3660 17604
rect 6828 17620 6880 17672
rect 9404 17620 9456 17672
rect 6000 17552 6052 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2044 17527 2096 17536
rect 2044 17493 2053 17527
rect 2053 17493 2087 17527
rect 2087 17493 2096 17527
rect 2044 17484 2096 17493
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2596 17323 2648 17332
rect 2596 17289 2605 17323
rect 2605 17289 2639 17323
rect 2639 17289 2648 17323
rect 2596 17280 2648 17289
rect 3608 17323 3660 17332
rect 3608 17289 3617 17323
rect 3617 17289 3651 17323
rect 3651 17289 3660 17323
rect 3608 17280 3660 17289
rect 7288 17323 7340 17332
rect 7288 17289 7297 17323
rect 7297 17289 7331 17323
rect 7331 17289 7340 17323
rect 7288 17280 7340 17289
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 4160 17076 4212 17128
rect 4252 17008 4304 17060
rect 5908 17144 5960 17196
rect 12164 17144 12216 17196
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 6000 16736 6052 16788
rect 12072 16668 12124 16720
rect 20720 16600 20772 16652
rect 21180 16600 21232 16652
rect 2412 16532 2464 16584
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 7196 16575 7248 16584
rect 7196 16541 7205 16575
rect 7205 16541 7239 16575
rect 7239 16541 7248 16575
rect 7196 16532 7248 16541
rect 8484 16532 8536 16584
rect 6920 16464 6972 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 6828 16396 6880 16448
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 8576 16396 8628 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 1676 16192 1728 16244
rect 1952 16099 2004 16108
rect 1952 16065 1961 16099
rect 1961 16065 1995 16099
rect 1995 16065 2004 16099
rect 1952 16056 2004 16065
rect 5172 16056 5224 16108
rect 2320 15988 2372 16040
rect 7656 15988 7708 16040
rect 2136 15963 2188 15972
rect 2136 15929 2145 15963
rect 2145 15929 2179 15963
rect 2179 15929 2188 15963
rect 2136 15920 2188 15929
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 5908 15648 5960 15700
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 12256 15512 12308 15564
rect 3792 15376 3844 15428
rect 7472 15444 7524 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 6000 15376 6052 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 9312 15308 9364 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 1676 15104 1728 15156
rect 2320 15104 2372 15156
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 3792 15147 3844 15156
rect 3792 15113 3801 15147
rect 3801 15113 3835 15147
rect 3835 15113 3844 15147
rect 3792 15104 3844 15113
rect 4160 15104 4212 15156
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 2412 14900 2464 14952
rect 4896 14968 4948 15020
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 5172 14832 5224 14884
rect 15384 15036 15436 15088
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 7380 14943 7432 14952
rect 5908 14900 5960 14909
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 7012 14832 7064 14884
rect 15568 14900 15620 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 2136 14560 2188 14612
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 9680 14560 9732 14612
rect 11704 14560 11756 14612
rect 4804 14492 4856 14544
rect 13268 14560 13320 14612
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 7104 14356 7156 14408
rect 10876 14424 10928 14476
rect 10508 14356 10560 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2136 14263 2188 14272
rect 2136 14229 2145 14263
rect 2145 14229 2179 14263
rect 2179 14229 2188 14263
rect 2136 14220 2188 14229
rect 2596 14220 2648 14272
rect 3976 14288 4028 14340
rect 4068 14220 4120 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 8300 14288 8352 14340
rect 4252 14220 4304 14229
rect 9680 14263 9732 14272
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 10324 14263 10376 14272
rect 9772 14220 9824 14229
rect 10324 14229 10333 14263
rect 10333 14229 10367 14263
rect 10367 14229 10376 14263
rect 10324 14220 10376 14229
rect 10784 14220 10836 14272
rect 12900 14220 12952 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 7380 14016 7432 14068
rect 8300 14059 8352 14068
rect 2780 13948 2832 14000
rect 6276 13948 6328 14000
rect 8300 14025 8309 14059
rect 8309 14025 8343 14059
rect 8343 14025 8352 14059
rect 8300 14016 8352 14025
rect 9404 14059 9456 14068
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 10324 14016 10376 14068
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10784 14059 10836 14068
rect 10416 14016 10468 14025
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 8116 13948 8168 14000
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3332 13880 3384 13932
rect 5264 13923 5316 13932
rect 3240 13812 3292 13864
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 5356 13855 5408 13864
rect 1860 13744 1912 13796
rect 3148 13744 3200 13796
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 5908 13812 5960 13864
rect 12900 14059 12952 14068
rect 12900 14025 12909 14059
rect 12909 14025 12943 14059
rect 12943 14025 12952 14059
rect 12900 14016 12952 14025
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 10968 13812 11020 13864
rect 8576 13744 8628 13796
rect 10140 13744 10192 13796
rect 4896 13676 4948 13728
rect 11152 13812 11204 13864
rect 11980 13744 12032 13796
rect 12348 13812 12400 13864
rect 12992 13676 13044 13728
rect 15660 13676 15712 13728
rect 18972 13676 19024 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 3240 13515 3292 13524
rect 2780 13472 2832 13481
rect 3240 13481 3249 13515
rect 3249 13481 3283 13515
rect 3283 13481 3292 13515
rect 3240 13472 3292 13481
rect 4252 13472 4304 13524
rect 7196 13472 7248 13524
rect 8576 13472 8628 13524
rect 11796 13472 11848 13524
rect 12072 13515 12124 13524
rect 12072 13481 12081 13515
rect 12081 13481 12115 13515
rect 12115 13481 12124 13515
rect 12072 13472 12124 13481
rect 2596 13336 2648 13388
rect 7840 13404 7892 13456
rect 3148 13336 3200 13388
rect 2964 13311 3016 13320
rect 1768 13132 1820 13184
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4436 13268 4488 13320
rect 4896 13336 4948 13388
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 6828 13336 6880 13388
rect 8208 13336 8260 13388
rect 5632 13268 5684 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 11060 13404 11112 13456
rect 11888 13404 11940 13456
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 17868 13336 17920 13388
rect 19708 13268 19760 13320
rect 3332 13200 3384 13252
rect 5356 13200 5408 13252
rect 2320 13132 2372 13184
rect 2412 13132 2464 13184
rect 4988 13132 5040 13184
rect 5448 13132 5500 13184
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 11704 13200 11756 13252
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 13084 13175 13136 13184
rect 12532 13132 12584 13141
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 20720 13132 20772 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 1676 12928 1728 12980
rect 7840 12971 7892 12980
rect 2872 12860 2924 12912
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 6828 12860 6880 12912
rect 4344 12792 4396 12844
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 6644 12767 6696 12776
rect 20 12656 72 12708
rect 4896 12656 4948 12708
rect 3332 12588 3384 12640
rect 4804 12588 4856 12640
rect 5632 12656 5684 12708
rect 6644 12733 6653 12767
rect 6653 12733 6687 12767
rect 6687 12733 6696 12767
rect 6644 12724 6696 12733
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 6920 12656 6972 12708
rect 8024 12724 8076 12776
rect 8208 12656 8260 12708
rect 11060 12928 11112 12980
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 13084 12928 13136 12980
rect 12072 12860 12124 12912
rect 9128 12792 9180 12844
rect 9680 12724 9732 12776
rect 10416 12724 10468 12776
rect 16764 12724 16816 12776
rect 21548 12656 21600 12708
rect 18420 12588 18472 12640
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 5724 12384 5776 12436
rect 6552 12384 6604 12436
rect 2504 12316 2556 12368
rect 8024 12384 8076 12436
rect 8484 12384 8536 12436
rect 11796 12384 11848 12436
rect 13176 12384 13228 12436
rect 13820 12384 13872 12436
rect 19064 12384 19116 12436
rect 2596 12248 2648 12300
rect 2780 12248 2832 12300
rect 3700 12248 3752 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 2872 12180 2924 12232
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 2780 12112 2832 12164
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 9956 12316 10008 12368
rect 8116 12248 8168 12300
rect 9588 12248 9640 12300
rect 11060 12248 11112 12300
rect 6920 12180 6972 12232
rect 7104 12180 7156 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 7748 12112 7800 12164
rect 8024 12112 8076 12164
rect 11704 12180 11756 12232
rect 20536 12223 20588 12232
rect 9864 12112 9916 12164
rect 12256 12112 12308 12164
rect 2136 12087 2188 12096
rect 2136 12053 2145 12087
rect 2145 12053 2179 12087
rect 2179 12053 2188 12087
rect 2136 12044 2188 12053
rect 2688 12044 2740 12096
rect 4988 12044 5040 12096
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 5540 12044 5592 12096
rect 5908 12044 5960 12096
rect 6552 12044 6604 12096
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7380 12044 7432 12096
rect 7932 12044 7984 12096
rect 9128 12044 9180 12096
rect 10600 12044 10652 12096
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 12164 12044 12216 12096
rect 14372 12112 14424 12164
rect 16764 12155 16816 12164
rect 16764 12121 16804 12155
rect 16804 12121 16816 12155
rect 16764 12112 16816 12121
rect 17316 12112 17368 12164
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 14280 12044 14332 12096
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 21456 12180 21508 12232
rect 20720 12112 20772 12164
rect 18328 12044 18380 12096
rect 21088 12044 21140 12096
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2136 11840 2188 11892
rect 2964 11840 3016 11892
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5448 11883 5500 11892
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 6000 11840 6052 11892
rect 6644 11840 6696 11892
rect 7380 11840 7432 11892
rect 7472 11840 7524 11892
rect 9220 11883 9272 11892
rect 9220 11849 9229 11883
rect 9229 11849 9263 11883
rect 9263 11849 9272 11883
rect 9220 11840 9272 11849
rect 2596 11772 2648 11824
rect 1492 11704 1544 11756
rect 2964 11704 3016 11756
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 2596 11636 2648 11645
rect 2780 11636 2832 11688
rect 5356 11815 5408 11824
rect 4620 11704 4672 11756
rect 5356 11781 5365 11815
rect 5365 11781 5399 11815
rect 5399 11781 5408 11815
rect 5356 11772 5408 11781
rect 9864 11840 9916 11892
rect 9956 11840 10008 11892
rect 15568 11883 15620 11892
rect 5908 11704 5960 11756
rect 8668 11704 8720 11756
rect 5632 11679 5684 11688
rect 3792 11568 3844 11620
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 7104 11636 7156 11688
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 13360 11772 13412 11824
rect 9128 11704 9180 11713
rect 11244 11704 11296 11756
rect 11704 11704 11756 11756
rect 13176 11704 13228 11756
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 2044 11500 2096 11552
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4160 11500 4212 11552
rect 7840 11500 7892 11552
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 18972 11840 19024 11892
rect 13728 11704 13780 11756
rect 14280 11704 14332 11756
rect 18328 11772 18380 11824
rect 20812 11772 20864 11824
rect 16488 11636 16540 11688
rect 12256 11500 12308 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 13820 11500 13872 11552
rect 18236 11704 18288 11756
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 18328 11636 18380 11645
rect 18144 11500 18196 11552
rect 19800 11500 19852 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 2964 11296 3016 11348
rect 4436 11296 4488 11348
rect 12164 11296 12216 11348
rect 3056 11228 3108 11280
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 2596 11160 2648 11212
rect 2780 11160 2832 11212
rect 5816 11160 5868 11212
rect 2228 11092 2280 11144
rect 8208 11228 8260 11280
rect 10600 11228 10652 11280
rect 6644 11160 6696 11212
rect 8024 11160 8076 11212
rect 8668 11160 8720 11212
rect 3424 11024 3476 11076
rect 4804 11024 4856 11076
rect 9128 11092 9180 11144
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 10968 11135 11020 11144
rect 10968 11101 11002 11135
rect 11002 11101 11020 11135
rect 15476 11296 15528 11348
rect 16488 11296 16540 11348
rect 19064 11296 19116 11348
rect 20812 11296 20864 11348
rect 12716 11228 12768 11280
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 21364 11296 21416 11348
rect 10968 11092 11020 11101
rect 13176 11092 13228 11144
rect 7104 11024 7156 11076
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 2780 10999 2832 11008
rect 2780 10965 2789 10999
rect 2789 10965 2823 10999
rect 2823 10965 2832 10999
rect 4896 10999 4948 11008
rect 2780 10956 2832 10965
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6552 10999 6604 11008
rect 6000 10956 6052 10965
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 6920 10956 6972 11008
rect 8208 10956 8260 11008
rect 12164 11024 12216 11076
rect 13360 11024 13412 11076
rect 15568 11135 15620 11144
rect 15568 11101 15586 11135
rect 15586 11101 15620 11135
rect 15568 11092 15620 11101
rect 18328 11092 18380 11144
rect 16396 11067 16448 11076
rect 16396 11033 16430 11067
rect 16430 11033 16448 11067
rect 16396 11024 16448 11033
rect 17040 11024 17092 11076
rect 18972 11024 19024 11076
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 1492 10752 1544 10804
rect 2136 10752 2188 10804
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 3148 10752 3200 10804
rect 3976 10752 4028 10804
rect 4896 10752 4948 10804
rect 2780 10684 2832 10736
rect 2044 10616 2096 10668
rect 2596 10591 2648 10600
rect 2596 10557 2605 10591
rect 2605 10557 2639 10591
rect 2639 10557 2648 10591
rect 2596 10548 2648 10557
rect 6644 10684 6696 10736
rect 11152 10752 11204 10804
rect 8944 10727 8996 10736
rect 8944 10693 8953 10727
rect 8953 10693 8987 10727
rect 8987 10693 8996 10727
rect 8944 10684 8996 10693
rect 15660 10752 15712 10804
rect 18236 10752 18288 10804
rect 3976 10616 4028 10668
rect 4068 10616 4120 10668
rect 5724 10616 5776 10668
rect 6920 10616 6972 10668
rect 9312 10616 9364 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 5448 10548 5500 10600
rect 6920 10480 6972 10532
rect 2412 10412 2464 10464
rect 5356 10412 5408 10464
rect 6828 10412 6880 10464
rect 8300 10412 8352 10464
rect 15476 10616 15528 10668
rect 15844 10659 15896 10668
rect 15844 10625 15862 10659
rect 15862 10625 15896 10659
rect 15844 10616 15896 10625
rect 17776 10659 17828 10668
rect 17776 10625 17794 10659
rect 17794 10625 17828 10659
rect 17776 10616 17828 10625
rect 19616 10616 19668 10668
rect 19800 10616 19852 10668
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 16304 10548 16356 10600
rect 9864 10412 9916 10464
rect 10232 10412 10284 10464
rect 12992 10412 13044 10464
rect 13084 10455 13136 10464
rect 13084 10421 13093 10455
rect 13093 10421 13127 10455
rect 13127 10421 13136 10455
rect 13084 10412 13136 10421
rect 13452 10412 13504 10464
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 16396 10412 16448 10464
rect 19064 10412 19116 10464
rect 19984 10455 20036 10464
rect 19984 10421 19993 10455
rect 19993 10421 20027 10455
rect 20027 10421 20036 10455
rect 19984 10412 20036 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1676 10208 1728 10260
rect 4068 10208 4120 10260
rect 6000 10208 6052 10260
rect 7288 10208 7340 10260
rect 2136 10140 2188 10192
rect 2320 10140 2372 10192
rect 3516 10140 3568 10192
rect 4160 10140 4212 10192
rect 5816 10140 5868 10192
rect 11888 10208 11940 10260
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 12992 10140 13044 10192
rect 19064 10208 19116 10260
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 5172 10072 5224 10124
rect 8024 10072 8076 10124
rect 8208 10072 8260 10124
rect 9680 10072 9732 10124
rect 21364 10251 21416 10260
rect 21364 10217 21373 10251
rect 21373 10217 21407 10251
rect 21407 10217 21416 10251
rect 21364 10208 21416 10217
rect 20720 10140 20772 10192
rect 1308 10004 1360 10056
rect 1492 10004 1544 10056
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 4068 10004 4120 10056
rect 5724 10004 5776 10056
rect 1952 9936 2004 9988
rect 4804 9979 4856 9988
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 2504 9868 2556 9877
rect 3056 9868 3108 9920
rect 4804 9945 4813 9979
rect 4813 9945 4847 9979
rect 4847 9945 4856 9979
rect 4804 9936 4856 9945
rect 5540 9936 5592 9988
rect 10692 10004 10744 10056
rect 12256 10004 12308 10056
rect 18420 10047 18472 10056
rect 18420 10013 18438 10047
rect 18438 10013 18472 10047
rect 18420 10004 18472 10013
rect 7104 9936 7156 9988
rect 11152 9936 11204 9988
rect 11704 9936 11756 9988
rect 16672 9979 16724 9988
rect 16672 9945 16681 9979
rect 16681 9945 16715 9979
rect 16715 9945 16724 9979
rect 16672 9936 16724 9945
rect 19248 9936 19300 9988
rect 19340 9936 19392 9988
rect 19708 9936 19760 9988
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 4988 9868 5040 9920
rect 5908 9868 5960 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 7564 9868 7616 9877
rect 7656 9868 7708 9920
rect 7932 9868 7984 9920
rect 8392 9868 8444 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9956 9911 10008 9920
rect 9404 9868 9456 9877
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 9956 9868 10008 9877
rect 12256 9868 12308 9920
rect 12808 9868 12860 9920
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 20168 9868 20220 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 1492 9664 1544 9716
rect 7564 9664 7616 9716
rect 9956 9664 10008 9716
rect 11060 9664 11112 9716
rect 19340 9707 19392 9716
rect 19340 9673 19349 9707
rect 19349 9673 19383 9707
rect 19383 9673 19392 9707
rect 19340 9664 19392 9673
rect 2044 9596 2096 9648
rect 2504 9596 2556 9648
rect 3148 9596 3200 9648
rect 4068 9596 4120 9648
rect 6920 9596 6972 9648
rect 8392 9639 8444 9648
rect 8392 9605 8401 9639
rect 8401 9605 8435 9639
rect 8435 9605 8444 9639
rect 8392 9596 8444 9605
rect 9864 9639 9916 9648
rect 9864 9605 9873 9639
rect 9873 9605 9907 9639
rect 9907 9605 9916 9639
rect 9864 9596 9916 9605
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 3240 9528 3292 9580
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5540 9528 5592 9580
rect 7656 9528 7708 9580
rect 2780 9460 2832 9512
rect 2872 9460 2924 9512
rect 3148 9460 3200 9512
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4160 9460 4212 9512
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 6920 9503 6972 9512
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 3332 9392 3384 9444
rect 5264 9392 5316 9444
rect 4528 9324 4580 9376
rect 4712 9324 4764 9376
rect 4988 9324 5040 9376
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 12440 9596 12492 9648
rect 10600 9528 10652 9580
rect 12164 9528 12216 9580
rect 14740 9596 14792 9648
rect 15568 9639 15620 9648
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 16304 9639 16356 9648
rect 15568 9596 15620 9605
rect 16304 9605 16313 9639
rect 16313 9605 16347 9639
rect 16347 9605 16356 9639
rect 16304 9596 16356 9605
rect 19248 9596 19300 9648
rect 20904 9664 20956 9716
rect 21364 9707 21416 9716
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 19984 9596 20036 9648
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 18144 9571 18196 9580
rect 18144 9537 18162 9571
rect 18162 9537 18196 9571
rect 18420 9571 18472 9580
rect 18144 9528 18196 9537
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 7012 9392 7064 9444
rect 10876 9503 10928 9512
rect 7564 9324 7616 9376
rect 9128 9324 9180 9376
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 11244 9324 11296 9376
rect 13176 9392 13228 9444
rect 17040 9435 17092 9444
rect 12624 9324 12676 9376
rect 15752 9324 15804 9376
rect 17040 9401 17049 9435
rect 17049 9401 17083 9435
rect 17083 9401 17092 9435
rect 17040 9392 17092 9401
rect 19524 9324 19576 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3976 9120 4028 9172
rect 6920 9120 6972 9172
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 7932 9052 7984 9104
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2596 8916 2648 8968
rect 4436 8916 4488 8968
rect 7656 8984 7708 9036
rect 8668 8916 8720 8968
rect 3332 8848 3384 8900
rect 6000 8848 6052 8900
rect 6736 8848 6788 8900
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 2320 8780 2372 8832
rect 2504 8780 2556 8832
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 3884 8780 3936 8832
rect 4436 8780 4488 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 5632 8780 5684 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 7564 8780 7616 8832
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8760 8780 8812 8832
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 10508 8916 10560 8968
rect 11152 8959 11204 8968
rect 10600 8780 10652 8832
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11336 9120 11388 9172
rect 11796 9120 11848 9172
rect 15936 9163 15988 9172
rect 15936 9129 15945 9163
rect 15945 9129 15979 9163
rect 15979 9129 15988 9163
rect 15936 9120 15988 9129
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 18420 9120 18472 9172
rect 19708 9163 19760 9172
rect 19708 9129 19717 9163
rect 19717 9129 19751 9163
rect 19751 9129 19760 9163
rect 19708 9120 19760 9129
rect 21364 8984 21416 9036
rect 12808 8959 12860 8968
rect 12072 8848 12124 8900
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 13820 8916 13872 8968
rect 20812 8959 20864 8968
rect 20812 8925 20830 8959
rect 20830 8925 20864 8959
rect 20812 8916 20864 8925
rect 12992 8848 13044 8900
rect 11796 8780 11848 8832
rect 14648 8848 14700 8900
rect 17960 8848 18012 8900
rect 14280 8780 14332 8832
rect 15752 8780 15804 8832
rect 20628 8780 20680 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 8392 8576 8444 8628
rect 8484 8576 8536 8628
rect 9496 8576 9548 8628
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 13452 8576 13504 8628
rect 1860 8508 1912 8560
rect 3884 8508 3936 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 1676 8372 1728 8424
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 4344 8415 4396 8424
rect 4068 8304 4120 8356
rect 4344 8381 4353 8415
rect 4353 8381 4387 8415
rect 4387 8381 4396 8415
rect 4344 8372 4396 8381
rect 4528 8508 4580 8560
rect 5172 8440 5224 8492
rect 10968 8508 11020 8560
rect 11888 8508 11940 8560
rect 8668 8440 8720 8492
rect 13176 8508 13228 8560
rect 15200 8576 15252 8628
rect 15568 8576 15620 8628
rect 15936 8576 15988 8628
rect 12992 8440 13044 8492
rect 13728 8440 13780 8492
rect 5632 8372 5684 8424
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8300 8372 8352 8424
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9864 8415 9916 8424
rect 5724 8304 5776 8356
rect 5816 8304 5868 8356
rect 6920 8304 6972 8356
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 11888 8372 11940 8424
rect 15200 8440 15252 8492
rect 15292 8372 15344 8424
rect 17868 8576 17920 8628
rect 17592 8508 17644 8560
rect 21180 8576 21232 8628
rect 18420 8440 18472 8492
rect 11796 8304 11848 8356
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 7472 8236 7524 8288
rect 12072 8304 12124 8356
rect 19524 8304 19576 8356
rect 12164 8236 12216 8288
rect 15844 8236 15896 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1400 8032 1452 8084
rect 4252 8032 4304 8084
rect 7564 8032 7616 8084
rect 1400 7871 1452 7880
rect 1400 7837 1433 7871
rect 1433 7837 1452 7871
rect 1860 7871 1912 7880
rect 1400 7828 1452 7837
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 5172 7896 5224 7948
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 5540 7896 5592 7948
rect 8576 8032 8628 8084
rect 9864 8032 9916 8084
rect 8300 7964 8352 8016
rect 2688 7828 2740 7880
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 3332 7828 3384 7880
rect 4712 7828 4764 7880
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 7288 7828 7340 7880
rect 1768 7692 1820 7744
rect 6828 7760 6880 7812
rect 9772 7828 9824 7880
rect 8116 7760 8168 7812
rect 11244 7896 11296 7948
rect 11704 7896 11756 7948
rect 15384 8032 15436 8084
rect 17316 8075 17368 8084
rect 15844 7964 15896 8016
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 12808 7828 12860 7880
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 17684 8032 17736 8084
rect 19616 8032 19668 8084
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 18512 8007 18564 8016
rect 18512 7973 18521 8007
rect 18521 7973 18555 8007
rect 18555 7973 18564 8007
rect 18512 7964 18564 7973
rect 21272 7964 21324 8016
rect 18420 7828 18472 7880
rect 2964 7692 3016 7744
rect 3976 7692 4028 7744
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 12164 7692 12216 7744
rect 12624 7760 12676 7812
rect 12900 7760 12952 7812
rect 14372 7760 14424 7812
rect 16304 7760 16356 7812
rect 19616 7760 19668 7812
rect 15844 7692 15896 7744
rect 19708 7692 19760 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 2596 7488 2648 7540
rect 4252 7488 4304 7540
rect 4344 7488 4396 7540
rect 4896 7488 4948 7540
rect 5264 7488 5316 7540
rect 5540 7488 5592 7540
rect 7196 7488 7248 7540
rect 8208 7488 8260 7540
rect 4988 7420 5040 7472
rect 5448 7420 5500 7472
rect 7380 7420 7432 7472
rect 8024 7420 8076 7472
rect 10692 7488 10744 7540
rect 11704 7488 11756 7540
rect 12440 7488 12492 7540
rect 15292 7531 15344 7540
rect 9680 7420 9732 7472
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 15936 7488 15988 7540
rect 16396 7488 16448 7540
rect 17684 7488 17736 7540
rect 17960 7488 18012 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1584 7352 1636 7404
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 2412 7352 2464 7404
rect 3240 7352 3292 7404
rect 4252 7352 4304 7404
rect 6368 7352 6420 7404
rect 8300 7395 8352 7404
rect 4804 7327 4856 7336
rect 1676 7216 1728 7268
rect 1860 7216 1912 7268
rect 2964 7259 3016 7268
rect 2964 7225 2973 7259
rect 2973 7225 3007 7259
rect 3007 7225 3016 7259
rect 2964 7216 3016 7225
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 7012 7284 7064 7336
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 12072 7352 12124 7404
rect 12624 7395 12676 7404
rect 12624 7361 12642 7395
rect 12642 7361 12676 7395
rect 12624 7352 12676 7361
rect 12808 7352 12860 7404
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 9404 7284 9456 7293
rect 10140 7284 10192 7336
rect 17684 7352 17736 7404
rect 19524 7420 19576 7472
rect 5172 7216 5224 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 7656 7148 7708 7200
rect 8208 7148 8260 7200
rect 10232 7191 10284 7200
rect 10232 7157 10241 7191
rect 10241 7157 10275 7191
rect 10275 7157 10284 7191
rect 10232 7148 10284 7157
rect 10416 7148 10468 7200
rect 13176 7216 13228 7268
rect 16212 7216 16264 7268
rect 21364 7488 21416 7540
rect 16764 7148 16816 7200
rect 19524 7148 19576 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2228 6944 2280 6996
rect 2688 6944 2740 6996
rect 4988 6944 5040 6996
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 2780 6808 2832 6860
rect 4160 6876 4212 6928
rect 4896 6876 4948 6928
rect 6828 6944 6880 6996
rect 8300 6944 8352 6996
rect 5632 6876 5684 6928
rect 16212 6944 16264 6996
rect 16396 6987 16448 6996
rect 16396 6953 16405 6987
rect 16405 6953 16439 6987
rect 16439 6953 16448 6987
rect 16396 6944 16448 6953
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3424 6740 3476 6792
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 6828 6851 6880 6860
rect 6828 6817 6837 6851
rect 6837 6817 6871 6851
rect 6871 6817 6880 6851
rect 6828 6808 6880 6817
rect 6368 6740 6420 6792
rect 8208 6808 8260 6860
rect 13176 6876 13228 6928
rect 7480 6779 7532 6788
rect 7480 6745 7489 6779
rect 7489 6745 7523 6779
rect 7523 6745 7532 6779
rect 7480 6736 7532 6745
rect 9404 6740 9456 6792
rect 11152 6808 11204 6860
rect 16028 6851 16080 6860
rect 16028 6817 16037 6851
rect 16037 6817 16071 6851
rect 16071 6817 16080 6851
rect 19524 6944 19576 6996
rect 21364 6987 21416 6996
rect 21364 6953 21373 6987
rect 21373 6953 21407 6987
rect 21407 6953 21416 6987
rect 21364 6944 21416 6953
rect 16028 6808 16080 6817
rect 18144 6851 18196 6860
rect 18144 6817 18153 6851
rect 18153 6817 18187 6851
rect 18187 6817 18196 6851
rect 18144 6808 18196 6817
rect 20996 6851 21048 6860
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 11704 6740 11756 6792
rect 4068 6604 4120 6656
rect 5908 6672 5960 6724
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 5172 6604 5224 6656
rect 5724 6604 5776 6656
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 7288 6647 7340 6656
rect 6736 6604 6788 6613
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 7380 6604 7432 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 9036 6604 9088 6656
rect 9956 6647 10008 6656
rect 9956 6613 9965 6647
rect 9965 6613 9999 6647
rect 9999 6613 10008 6647
rect 9956 6604 10008 6613
rect 10968 6604 11020 6656
rect 15200 6672 15252 6724
rect 15752 6715 15804 6724
rect 15752 6681 15770 6715
rect 15770 6681 15804 6715
rect 15752 6672 15804 6681
rect 14648 6647 14700 6656
rect 14648 6613 14657 6647
rect 14657 6613 14691 6647
rect 14691 6613 14700 6647
rect 14648 6604 14700 6613
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 17316 6604 17368 6656
rect 18052 6672 18104 6724
rect 19708 6672 19760 6724
rect 18328 6604 18380 6656
rect 18972 6604 19024 6656
rect 19616 6604 19668 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 5540 6400 5592 6452
rect 5724 6400 5776 6452
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 6736 6443 6788 6452
rect 6736 6409 6745 6443
rect 6745 6409 6779 6443
rect 6779 6409 6788 6443
rect 6736 6400 6788 6409
rect 8116 6400 8168 6452
rect 9036 6443 9088 6452
rect 8668 6375 8720 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 1768 6196 1820 6248
rect 2872 6196 2924 6248
rect 3332 6264 3384 6316
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4528 6264 4580 6316
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 8668 6341 8677 6375
rect 8677 6341 8711 6375
rect 8711 6341 8720 6375
rect 8668 6332 8720 6341
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 11152 6400 11204 6452
rect 11704 6400 11756 6452
rect 13176 6400 13228 6452
rect 9312 6332 9364 6384
rect 9956 6332 10008 6384
rect 12808 6332 12860 6384
rect 10232 6264 10284 6316
rect 11704 6264 11756 6316
rect 12164 6264 12216 6316
rect 13176 6264 13228 6316
rect 13360 6264 13412 6316
rect 14832 6307 14884 6316
rect 14832 6273 14850 6307
rect 14850 6273 14884 6307
rect 14832 6264 14884 6273
rect 15200 6264 15252 6316
rect 16028 6400 16080 6452
rect 3056 6196 3108 6248
rect 5264 6196 5316 6248
rect 2044 6128 2096 6180
rect 5632 6128 5684 6180
rect 5908 6196 5960 6248
rect 7380 6239 7432 6248
rect 6460 6128 6512 6180
rect 6552 6128 6604 6180
rect 7012 6128 7064 6180
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 9312 6239 9364 6248
rect 7564 6128 7616 6180
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 13636 6196 13688 6248
rect 18144 6400 18196 6452
rect 18972 6332 19024 6384
rect 16948 6307 17000 6316
rect 16948 6273 16982 6307
rect 16982 6273 17000 6307
rect 16948 6264 17000 6273
rect 17408 6264 17460 6316
rect 19248 6400 19300 6452
rect 20444 6400 20496 6452
rect 21088 6264 21140 6316
rect 1676 6060 1728 6112
rect 3240 6060 3292 6112
rect 4068 6060 4120 6112
rect 4896 6060 4948 6112
rect 5540 6060 5592 6112
rect 6736 6060 6788 6112
rect 9496 6060 9548 6112
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 11796 6060 11848 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 13728 6103 13780 6112
rect 11888 6060 11940 6069
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 13728 6060 13780 6069
rect 13820 6060 13872 6112
rect 17592 6060 17644 6112
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 2320 5856 2372 5908
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 2596 5788 2648 5840
rect 3240 5788 3292 5840
rect 4528 5720 4580 5772
rect 6828 5856 6880 5908
rect 8760 5856 8812 5908
rect 8300 5788 8352 5840
rect 6460 5720 6512 5772
rect 9496 5856 9548 5908
rect 9864 5856 9916 5908
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 13360 5899 13412 5908
rect 13360 5865 13369 5899
rect 13369 5865 13403 5899
rect 13403 5865 13412 5899
rect 13360 5856 13412 5865
rect 13636 5856 13688 5908
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 3516 5652 3568 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4068 5652 4120 5704
rect 7840 5652 7892 5704
rect 14372 5788 14424 5840
rect 16028 5856 16080 5908
rect 19708 5856 19760 5908
rect 19800 5856 19852 5908
rect 20996 5788 21048 5840
rect 9036 5720 9088 5772
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 1676 5627 1728 5636
rect 1676 5593 1685 5627
rect 1685 5593 1719 5627
rect 1719 5593 1728 5627
rect 1676 5584 1728 5593
rect 3240 5584 3292 5636
rect 2412 5516 2464 5568
rect 2964 5516 3016 5568
rect 3608 5516 3660 5568
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 5172 5516 5224 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 5724 5516 5776 5568
rect 7932 5584 7984 5636
rect 13360 5720 13412 5772
rect 14464 5720 14516 5772
rect 16028 5720 16080 5772
rect 13728 5652 13780 5704
rect 17592 5652 17644 5704
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 10968 5516 11020 5568
rect 14280 5584 14332 5636
rect 15568 5584 15620 5636
rect 15752 5584 15804 5636
rect 17960 5584 18012 5636
rect 19432 5652 19484 5704
rect 20076 5584 20128 5636
rect 20444 5627 20496 5636
rect 20444 5593 20462 5627
rect 20462 5593 20496 5627
rect 20444 5584 20496 5593
rect 13820 5516 13872 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14372 5516 14424 5568
rect 18236 5516 18288 5568
rect 19248 5516 19300 5568
rect 20720 5516 20772 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2596 5355 2648 5364
rect 2596 5321 2605 5355
rect 2605 5321 2639 5355
rect 2639 5321 2648 5355
rect 2596 5312 2648 5321
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 3516 5312 3568 5364
rect 4068 5312 4120 5364
rect 4804 5312 4856 5364
rect 5264 5312 5316 5364
rect 5908 5312 5960 5364
rect 6092 5312 6144 5364
rect 6552 5312 6604 5364
rect 3424 5244 3476 5296
rect 8116 5312 8168 5364
rect 9956 5312 10008 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 4712 5176 4764 5228
rect 4804 5176 4856 5228
rect 7932 5244 7984 5296
rect 5632 5176 5684 5228
rect 3148 5108 3200 5160
rect 3608 5108 3660 5160
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5908 5108 5960 5160
rect 8484 5176 8536 5228
rect 10048 5176 10100 5228
rect 5264 5040 5316 5092
rect 6736 5040 6788 5092
rect 8668 5108 8720 5160
rect 9128 5108 9180 5160
rect 11888 5312 11940 5364
rect 13360 5312 13412 5364
rect 16028 5312 16080 5364
rect 19432 5355 19484 5364
rect 19432 5321 19441 5355
rect 19441 5321 19475 5355
rect 19475 5321 19484 5355
rect 19432 5312 19484 5321
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 12624 5219 12676 5228
rect 12624 5185 12642 5219
rect 12642 5185 12676 5219
rect 12624 5176 12676 5185
rect 13360 5176 13412 5228
rect 14096 5176 14148 5228
rect 11704 5108 11756 5160
rect 17132 5244 17184 5296
rect 21180 5244 21232 5296
rect 18512 5176 18564 5228
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 20812 5219 20864 5228
rect 20812 5185 20830 5219
rect 20830 5185 20864 5219
rect 20812 5176 20864 5185
rect 20996 5176 21048 5228
rect 18052 5108 18104 5160
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 3976 4972 4028 5024
rect 4988 4972 5040 5024
rect 5632 4972 5684 5024
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7012 4972 7064 5024
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 8576 4972 8628 5024
rect 9404 4972 9456 5024
rect 9680 4972 9732 5024
rect 9956 4972 10008 5024
rect 11704 4972 11756 5024
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 15752 4972 15804 5024
rect 18512 5040 18564 5092
rect 18144 4972 18196 5024
rect 18604 4972 18656 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 2136 4632 2188 4684
rect 3148 4700 3200 4752
rect 4620 4768 4672 4820
rect 6828 4768 6880 4820
rect 1860 4564 1912 4616
rect 2964 4632 3016 4684
rect 2412 4564 2464 4616
rect 4436 4564 4488 4616
rect 5264 4564 5316 4616
rect 5540 4564 5592 4616
rect 6368 4632 6420 4684
rect 8392 4632 8444 4684
rect 6736 4564 6788 4616
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 12900 4768 12952 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 14280 4768 14332 4820
rect 12532 4700 12584 4752
rect 16304 4700 16356 4752
rect 10968 4632 11020 4684
rect 11152 4632 11204 4684
rect 10324 4564 10376 4616
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12808 4564 12860 4616
rect 5356 4496 5408 4548
rect 6092 4496 6144 4548
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 5080 4428 5132 4480
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 7380 4428 7432 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 8852 4428 8904 4480
rect 9496 4471 9548 4480
rect 9496 4437 9505 4471
rect 9505 4437 9539 4471
rect 9539 4437 9548 4471
rect 9496 4428 9548 4437
rect 9680 4428 9732 4480
rect 11060 4496 11112 4548
rect 11244 4496 11296 4548
rect 12348 4496 12400 4548
rect 13360 4496 13412 4548
rect 15752 4496 15804 4548
rect 16028 4564 16080 4616
rect 16948 4632 17000 4684
rect 18236 4768 18288 4820
rect 12440 4428 12492 4480
rect 13544 4428 13596 4480
rect 14372 4428 14424 4480
rect 18420 4496 18472 4548
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 17868 4428 17920 4480
rect 20996 4632 21048 4684
rect 21456 4564 21508 4616
rect 19708 4496 19760 4548
rect 21088 4471 21140 4480
rect 21088 4437 21097 4471
rect 21097 4437 21131 4471
rect 21131 4437 21140 4471
rect 21088 4428 21140 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 3424 4224 3476 4276
rect 4252 4224 4304 4276
rect 7564 4224 7616 4276
rect 1768 4088 1820 4140
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 3240 4088 3292 4140
rect 4344 4156 4396 4208
rect 4988 4156 5040 4208
rect 5632 4156 5684 4208
rect 6184 4156 6236 4208
rect 6920 4156 6972 4208
rect 3884 4088 3936 4140
rect 4160 4088 4212 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 5080 4088 5132 4140
rect 4068 4020 4120 4072
rect 6276 4088 6328 4140
rect 7196 4088 7248 4140
rect 7472 4088 7524 4140
rect 7656 4088 7708 4140
rect 12164 4224 12216 4276
rect 12348 4267 12400 4276
rect 12348 4233 12357 4267
rect 12357 4233 12391 4267
rect 12391 4233 12400 4267
rect 12348 4224 12400 4233
rect 12440 4224 12492 4276
rect 15108 4224 15160 4276
rect 9680 4156 9732 4208
rect 5908 4020 5960 4072
rect 6920 4063 6972 4072
rect 6920 4029 6929 4063
rect 6929 4029 6963 4063
rect 6963 4029 6972 4063
rect 6920 4020 6972 4029
rect 9128 4088 9180 4140
rect 9772 4088 9824 4140
rect 10692 4088 10744 4140
rect 10876 4088 10928 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 13360 4156 13412 4208
rect 3240 3952 3292 4004
rect 3608 3952 3660 4004
rect 3976 3995 4028 4004
rect 3976 3961 3985 3995
rect 3985 3961 4019 3995
rect 4019 3961 4028 3995
rect 3976 3952 4028 3961
rect 4436 3995 4488 4004
rect 4436 3961 4445 3995
rect 4445 3961 4479 3995
rect 4479 3961 4488 3995
rect 4436 3952 4488 3961
rect 4804 3952 4856 4004
rect 5172 3995 5224 4004
rect 5172 3961 5181 3995
rect 5181 3961 5215 3995
rect 5215 3961 5224 3995
rect 5172 3952 5224 3961
rect 5540 3952 5592 4004
rect 8852 4020 8904 4072
rect 3424 3884 3476 3936
rect 8024 3884 8076 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 9312 3952 9364 4004
rect 9956 3995 10008 4004
rect 9956 3961 9965 3995
rect 9965 3961 9999 3995
rect 9999 3961 10008 3995
rect 9956 3952 10008 3961
rect 12900 4020 12952 4072
rect 11060 3952 11112 4004
rect 11520 3952 11572 4004
rect 12808 3952 12860 4004
rect 10508 3884 10560 3936
rect 11336 3884 11388 3936
rect 11888 3884 11940 3936
rect 13268 4088 13320 4140
rect 14464 4156 14516 4208
rect 16856 4224 16908 4276
rect 17868 4224 17920 4276
rect 16028 4156 16080 4208
rect 20996 4156 21048 4208
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 17224 4088 17276 4140
rect 19432 4131 19484 4140
rect 19432 4097 19450 4131
rect 19450 4097 19484 4131
rect 19708 4131 19760 4140
rect 19432 4088 19484 4097
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 21272 4088 21324 4140
rect 16396 3884 16448 3936
rect 17960 3952 18012 4004
rect 17316 3884 17368 3936
rect 17776 3884 17828 3936
rect 18512 3884 18564 3936
rect 20 3748 72 3800
rect 940 3748 992 3800
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 4712 3680 4764 3732
rect 5540 3723 5592 3732
rect 5540 3689 5549 3723
rect 5549 3689 5583 3723
rect 5583 3689 5592 3723
rect 5540 3680 5592 3689
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 6276 3680 6328 3732
rect 6828 3680 6880 3732
rect 8300 3680 8352 3732
rect 8852 3680 8904 3732
rect 15936 3680 15988 3732
rect 16856 3680 16908 3732
rect 8944 3612 8996 3664
rect 9772 3612 9824 3664
rect 11336 3612 11388 3664
rect 14280 3612 14332 3664
rect 15568 3612 15620 3664
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 2964 3544 3016 3596
rect 940 3476 992 3528
rect 3240 3476 3292 3528
rect 3424 3476 3476 3528
rect 6092 3544 6144 3596
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 6552 3544 6604 3596
rect 7840 3544 7892 3596
rect 8116 3544 8168 3596
rect 8668 3544 8720 3596
rect 9404 3544 9456 3596
rect 9680 3544 9732 3596
rect 11152 3544 11204 3596
rect 16028 3544 16080 3596
rect 17132 3612 17184 3664
rect 18972 3680 19024 3732
rect 21088 3680 21140 3732
rect 18512 3544 18564 3596
rect 19616 3544 19668 3596
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 6644 3476 6696 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 8576 3519 8628 3528
rect 7564 3476 7616 3485
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 9036 3476 9088 3528
rect 5448 3408 5500 3460
rect 6092 3408 6144 3460
rect 6552 3408 6604 3460
rect 9588 3452 9640 3504
rect 10232 3476 10284 3528
rect 10692 3519 10744 3528
rect 10692 3485 10710 3519
rect 10710 3485 10744 3519
rect 10692 3476 10744 3485
rect 13544 3519 13596 3528
rect 10784 3408 10836 3460
rect 12532 3408 12584 3460
rect 5264 3340 5316 3392
rect 5908 3340 5960 3392
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 9496 3340 9548 3392
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 14648 3476 14700 3528
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 18420 3476 18472 3528
rect 20536 3476 20588 3528
rect 20996 3476 21048 3528
rect 15016 3408 15068 3460
rect 18144 3408 18196 3460
rect 18236 3408 18288 3460
rect 13820 3340 13872 3392
rect 16396 3340 16448 3392
rect 17500 3340 17552 3392
rect 19800 3408 19852 3460
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 6920 3136 6972 3188
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 8116 3179 8168 3188
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 8852 3136 8904 3188
rect 9312 3136 9364 3188
rect 9496 3179 9548 3188
rect 9496 3145 9505 3179
rect 9505 3145 9539 3179
rect 9539 3145 9548 3179
rect 9496 3136 9548 3145
rect 12348 3136 12400 3188
rect 2596 3068 2648 3120
rect 1492 3000 1544 3052
rect 3240 3000 3292 3052
rect 3700 3000 3752 3052
rect 7288 3068 7340 3120
rect 8944 3068 8996 3120
rect 2780 2932 2832 2984
rect 3148 2932 3200 2984
rect 3424 2932 3476 2984
rect 7104 3000 7156 3052
rect 8392 3043 8444 3052
rect 6736 2975 6788 2984
rect 6000 2907 6052 2916
rect 6000 2873 6009 2907
rect 6009 2873 6043 2907
rect 6043 2873 6052 2907
rect 6000 2864 6052 2873
rect 6736 2941 6745 2975
rect 6745 2941 6779 2975
rect 6779 2941 6788 2975
rect 6736 2932 6788 2941
rect 7840 2932 7892 2984
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 9220 3000 9272 3052
rect 9680 3000 9732 3052
rect 10508 3000 10560 3052
rect 10600 3000 10652 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 8668 2932 8720 2984
rect 9772 2932 9824 2984
rect 12900 3068 12952 3120
rect 16856 3136 16908 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 17868 3136 17920 3188
rect 21272 3136 21324 3188
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 15384 3043 15436 3052
rect 7564 2864 7616 2916
rect 8024 2864 8076 2916
rect 9220 2864 9272 2916
rect 7196 2796 7248 2848
rect 7656 2796 7708 2848
rect 7748 2796 7800 2848
rect 13360 2932 13412 2984
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 18328 3068 18380 3120
rect 14372 2932 14424 2984
rect 17040 2932 17092 2984
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 13268 2864 13320 2916
rect 17776 2932 17828 2984
rect 20812 3000 20864 3052
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 13452 2796 13504 2848
rect 14280 2796 14332 2848
rect 15292 2796 15344 2848
rect 15660 2796 15712 2848
rect 16948 2796 17000 2848
rect 19524 2796 19576 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 11152 2592 11204 2644
rect 2504 2524 2556 2576
rect 4804 2524 4856 2576
rect 6644 2524 6696 2576
rect 9220 2524 9272 2576
rect 2044 2388 2096 2440
rect 2320 2456 2372 2508
rect 2412 2456 2464 2508
rect 3976 2456 4028 2508
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 4804 2388 4856 2440
rect 7104 2456 7156 2508
rect 5540 2388 5592 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6828 2388 6880 2440
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 8484 2456 8536 2508
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 9864 2524 9916 2576
rect 11244 2524 11296 2576
rect 9588 2388 9640 2440
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 4068 2320 4120 2372
rect 4252 2320 4304 2372
rect 11796 2456 11848 2508
rect 16580 2592 16632 2644
rect 19340 2592 19392 2644
rect 13084 2524 13136 2576
rect 14556 2524 14608 2576
rect 16396 2524 16448 2576
rect 13820 2456 13872 2508
rect 11704 2388 11756 2440
rect 12808 2388 12860 2440
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 15108 2456 15160 2508
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 19708 2592 19760 2644
rect 20168 2592 20220 2644
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 15844 2388 15896 2440
rect 18328 2431 18380 2440
rect 1308 2252 1360 2304
rect 5908 2252 5960 2304
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 7472 2252 7524 2304
rect 7656 2295 7708 2304
rect 7656 2261 7665 2295
rect 7665 2261 7699 2295
rect 7699 2261 7708 2295
rect 7656 2252 7708 2261
rect 7932 2252 7984 2304
rect 9404 2252 9456 2304
rect 9680 2252 9732 2304
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 10692 2295 10744 2304
rect 10692 2261 10701 2295
rect 10701 2261 10735 2295
rect 10735 2261 10744 2295
rect 10692 2252 10744 2261
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 12808 2252 12860 2304
rect 13820 2320 13872 2372
rect 14372 2252 14424 2304
rect 15016 2320 15068 2372
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 19524 2388 19576 2440
rect 21456 2388 21508 2440
rect 18144 2320 18196 2372
rect 14924 2252 14976 2304
rect 16028 2252 16080 2304
rect 20720 2252 20772 2304
rect 20904 2252 20956 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 5540 2048 5592 2100
rect 8300 2048 8352 2100
rect 5448 1980 5500 2032
rect 13176 2048 13228 2100
rect 10048 1980 10100 2032
rect 17040 1980 17092 2032
rect 7472 1912 7524 1964
rect 15844 1912 15896 1964
rect 4068 1844 4120 1896
rect 4804 1844 4856 1896
rect 10416 1844 10468 1896
rect 10692 1844 10744 1896
rect 12440 1844 12492 1896
rect 5816 1776 5868 1828
rect 8668 1776 8720 1828
rect 7840 1708 7892 1760
rect 7104 1640 7156 1692
rect 7932 1640 7984 1692
rect 8208 1708 8260 1760
rect 14096 1776 14148 1828
rect 12072 1708 12124 1760
rect 15384 1708 15436 1760
rect 20720 1912 20772 1964
rect 11612 1572 11664 1624
rect 11796 1572 11848 1624
rect 18328 1640 18380 1692
rect 5724 1504 5776 1556
rect 6460 1504 6512 1556
rect 7656 1436 7708 1488
rect 12072 1436 12124 1488
rect 9680 1368 9732 1420
rect 9956 1368 10008 1420
<< metal2 >>
rect 2962 21312 3018 21321
rect 2962 21247 3018 21256
rect 2870 20904 2926 20913
rect 2870 20839 2926 20848
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2792 20505 2820 20538
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 1860 20392 1912 20398
rect 1860 20334 1912 20340
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1688 18970 1716 19790
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1490 18864 1546 18873
rect 1490 18799 1546 18808
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1688 17882 1716 18226
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1490 16759 1546 16768
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1688 16250 1716 17138
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15609 1532 15846
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1688 15162 1716 15438
rect 1490 15127 1546 15136
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13977 1532 14214
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13569 1532 13670
rect 1490 13560 1546 13569
rect 1490 13495 1546 13504
rect 1490 13152 1546 13161
rect 1490 13087 1546 13096
rect 1504 12986 1532 13087
rect 1688 12986 1716 14350
rect 1872 13802 1900 20334
rect 2042 20088 2098 20097
rect 2884 20058 2912 20839
rect 2976 20398 3004 21247
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 4448 20058 4476 20402
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 2042 20023 2044 20032
rect 2096 20023 2098 20032
rect 2872 20052 2924 20058
rect 2044 19994 2096 20000
rect 2872 19994 2924 20000
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 2240 19514 2268 19790
rect 5736 19514 5764 19790
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 1964 17814 1992 19314
rect 2042 19272 2098 19281
rect 2042 19207 2044 19216
rect 2096 19207 2098 19216
rect 2044 19178 2096 19184
rect 2240 18426 2268 19314
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3896 17882 3924 18702
rect 5920 17882 5948 18702
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 1952 17808 2004 17814
rect 1952 17750 2004 17756
rect 1952 17672 2004 17678
rect 2596 17672 2648 17678
rect 1952 17614 2004 17620
rect 2042 17640 2098 17649
rect 1964 17338 1992 17614
rect 2596 17614 2648 17620
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 2042 17575 2098 17584
rect 2056 17542 2084 17575
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2608 17338 2636 17614
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 3620 17338 3648 17546
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1964 15706 1992 16050
rect 2320 16040 2372 16046
rect 2134 16008 2190 16017
rect 2320 15982 2372 15988
rect 2134 15943 2136 15952
rect 2188 15943 2190 15952
rect 2136 15914 2188 15920
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2332 15162 2360 15982
rect 2424 15706 2452 16526
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3804 15162 3832 15370
rect 4172 15162 4200 17070
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4264 16794 4292 17002
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15706 5212 16050
rect 5920 15706 5948 17138
rect 6012 16794 6040 17546
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 2148 14618 2176 14962
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2134 14376 2190 14385
rect 1964 14074 1992 14350
rect 2134 14311 2190 14320
rect 2148 14278 2176 14311
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2424 14074 2452 14894
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 4816 14550 4844 14894
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2608 13938 2636 14214
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 2792 13530 2820 13942
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1398 12744 1454 12753
rect 20 12708 72 12714
rect 1398 12679 1454 12688
rect 20 12650 72 12656
rect 32 3806 60 12650
rect 1412 12238 1440 12679
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1214 11792 1270 11801
rect 1214 11727 1270 11736
rect 20 3800 72 3806
rect 940 3800 992 3806
rect 20 3742 72 3748
rect 938 3768 940 3777
rect 992 3768 994 3777
rect 938 3703 994 3712
rect 952 3534 980 3703
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 1228 2774 1256 11727
rect 1412 11354 1440 12174
rect 1504 11762 1532 12271
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1584 11552 1636 11558
rect 1490 11520 1546 11529
rect 1584 11494 1636 11500
rect 1490 11455 1546 11464
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1412 10418 1440 10911
rect 1504 10810 1532 11455
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1490 10704 1546 10713
rect 1490 10639 1546 10648
rect 1320 10390 1440 10418
rect 1320 10062 1348 10390
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1412 9586 1440 10231
rect 1504 10062 1532 10639
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9722 1532 9998
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1412 8974 1440 9007
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1412 8090 1440 8191
rect 1490 8120 1546 8129
rect 1400 8084 1452 8090
rect 1490 8055 1546 8064
rect 1400 8026 1452 8032
rect 1400 7880 1452 7886
rect 1398 7848 1400 7857
rect 1452 7848 1454 7857
rect 1398 7783 1454 7792
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 7041 1440 7346
rect 1398 7032 1454 7041
rect 1398 6967 1454 6976
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6633 1440 6734
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 6225 1440 6258
rect 1398 6216 1454 6225
rect 1398 6151 1454 6160
rect 1398 5400 1454 5409
rect 1398 5335 1454 5344
rect 1412 5234 1440 5335
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1504 3058 1532 8055
rect 1596 7410 1624 11494
rect 1674 10704 1730 10713
rect 1674 10639 1730 10648
rect 1688 10266 1716 10639
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1688 7274 1716 8366
rect 1780 7970 1808 13126
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11898 2176 12038
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1950 11248 2006 11257
rect 2056 11218 2084 11494
rect 1950 11183 1952 11192
rect 2004 11183 2006 11192
rect 2044 11212 2096 11218
rect 1952 11154 2004 11160
rect 2044 11154 2096 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2148 10810 2176 10950
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1872 9489 1900 9522
rect 1858 9480 1914 9489
rect 1858 9415 1914 9424
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 8673 1900 8910
rect 1858 8664 1914 8673
rect 1964 8634 1992 9930
rect 2056 9654 2084 10610
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9081 2084 9318
rect 2042 9072 2098 9081
rect 2042 9007 2098 9016
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1858 8599 1914 8608
rect 1952 8628 2004 8634
rect 1872 8566 1900 8599
rect 1952 8570 2004 8576
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 2056 8401 2084 8774
rect 2042 8392 2098 8401
rect 2042 8327 2098 8336
rect 2042 7984 2098 7993
rect 1780 7942 1992 7970
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7041 1624 7142
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1780 6361 1808 7686
rect 1872 7449 1900 7822
rect 1858 7440 1914 7449
rect 1858 7375 1914 7384
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1766 6352 1822 6361
rect 1766 6287 1822 6296
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1582 5672 1638 5681
rect 1688 5642 1716 6054
rect 1780 5710 1808 6190
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1582 5607 1638 5616
rect 1676 5636 1728 5642
rect 1596 5370 1624 5607
rect 1676 5578 1728 5584
rect 1872 5556 1900 7210
rect 1780 5528 1900 5556
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1780 4146 1808 5528
rect 1860 5024 1912 5030
rect 1858 4992 1860 5001
rect 1912 4992 1914 5001
rect 1858 4927 1914 4936
rect 1860 4616 1912 4622
rect 1858 4584 1860 4593
rect 1912 4584 1914 4593
rect 1858 4519 1914 4528
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1964 3602 1992 7942
rect 2042 7919 2098 7928
rect 2056 7546 2084 7919
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 2056 3641 2084 6122
rect 2148 4690 2176 10134
rect 2240 7002 2268 11086
rect 2332 10198 2360 13126
rect 2424 10810 2452 13126
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2332 9897 2360 9998
rect 2318 9888 2374 9897
rect 2318 9823 2374 9832
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8430 2360 8774
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2424 7410 2452 10406
rect 2516 10146 2544 12310
rect 2608 12306 2636 13330
rect 2884 12918 2912 13670
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2608 11830 2636 12242
rect 2792 12170 2820 12242
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2596 11688 2648 11694
rect 2594 11656 2596 11665
rect 2648 11656 2650 11665
rect 2594 11591 2650 11600
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 10606 2636 11154
rect 2596 10600 2648 10606
rect 2594 10568 2596 10577
rect 2648 10568 2650 10577
rect 2594 10503 2650 10512
rect 2516 10118 2636 10146
rect 2502 10024 2558 10033
rect 2502 9959 2558 9968
rect 2516 9926 2544 9959
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2516 8838 2544 9590
rect 2608 8974 2636 10118
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2700 7886 2728 12038
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 11218 2820 11630
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10742 2820 10950
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2884 9518 2912 12174
rect 2976 11898 3004 13262
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11354 3004 11698
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 3068 11286 3096 13874
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3160 13394 3188 13738
rect 3252 13530 3280 13806
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3344 13258 3372 13874
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12238 3372 12582
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 11937 3372 12174
rect 3330 11928 3386 11937
rect 3330 11863 3386 11872
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2962 10160 3018 10169
rect 2962 10095 3018 10104
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2792 7886 2820 9454
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8634 2912 8774
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2688 7880 2740 7886
rect 2502 7848 2558 7857
rect 2688 7822 2740 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2502 7783 2558 7792
rect 2516 7546 2544 7783
rect 2976 7750 3004 10095
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 8129 3096 9862
rect 3160 9654 3188 10746
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 9058 3188 9454
rect 3252 9178 3280 9522
rect 3344 9450 3372 11698
rect 3712 11558 3740 12242
rect 3882 12200 3938 12209
rect 3882 12135 3938 12144
rect 3790 11656 3846 11665
rect 3790 11591 3792 11600
rect 3844 11591 3846 11600
rect 3792 11562 3844 11568
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3160 9030 3280 9058
rect 3054 8120 3110 8129
rect 3054 8055 3110 8064
rect 3252 7868 3280 9030
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 7886 3372 8842
rect 3160 7840 3280 7868
rect 3332 7880 3384 7886
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2870 7576 2926 7585
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2596 7540 2648 7546
rect 2870 7511 2926 7520
rect 2596 7482 2648 7488
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2412 7404 2464 7410
rect 2608 7392 2636 7482
rect 2412 7346 2464 7352
rect 2516 7364 2636 7392
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2226 6896 2282 6905
rect 2226 6831 2228 6840
rect 2280 6831 2282 6840
rect 2228 6802 2280 6808
rect 2332 5914 2360 7346
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2318 5128 2374 5137
rect 2318 5063 2374 5072
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2226 4176 2282 4185
rect 2226 4111 2228 4120
rect 2280 4111 2282 4120
rect 2228 4082 2280 4088
rect 2042 3632 2098 3641
rect 1952 3596 2004 3602
rect 2042 3567 2098 3576
rect 1952 3538 2004 3544
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1228 2746 1348 2774
rect 1320 2310 1348 2746
rect 2332 2514 2360 5063
rect 2424 4622 2452 5510
rect 2516 5234 2544 7364
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2608 5370 2636 5782
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2516 2582 2544 5170
rect 2700 4978 2728 6938
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2792 6322 2820 6802
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2792 5817 2820 6258
rect 2884 6254 2912 7511
rect 2962 7304 3018 7313
rect 2962 7239 2964 7248
rect 3016 7239 3018 7248
rect 2964 7210 3016 7216
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2792 5001 2820 5199
rect 2608 4950 2728 4978
rect 2778 4992 2834 5001
rect 2608 3126 2636 4950
rect 2778 4927 2834 4936
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2778 3088 2834 3097
rect 2778 3023 2834 3032
rect 2792 2990 2820 3023
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2884 2836 2912 6190
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5370 3004 5510
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2962 4992 3018 5001
rect 2962 4927 3018 4936
rect 2976 4690 3004 4927
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2962 4584 3018 4593
rect 2962 4519 3018 4528
rect 2976 3602 3004 4519
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2792 2808 2912 2836
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 2056 800 2084 2382
rect 2424 800 2452 2450
rect 2792 800 2820 2808
rect 2976 2553 3004 3538
rect 3068 2774 3096 6190
rect 3160 5522 3188 7840
rect 3332 7822 3384 7828
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 6118 3280 7346
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6322 3372 7142
rect 3436 6798 3464 11018
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3528 9489 3556 10134
rect 3514 9480 3570 9489
rect 3514 9415 3570 9424
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3896 8838 3924 12135
rect 3988 10810 4016 14282
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4080 14074 4108 14214
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4264 13530 4292 14214
rect 4908 14074 4936 14962
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4908 13394 4936 13670
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4356 12442 4384 12786
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3988 10130 4016 10610
rect 4080 10266 4108 10610
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4172 10198 4200 11494
rect 4448 11354 4476 13262
rect 4908 12714 4936 13330
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4816 12306 4844 12582
rect 5000 12434 5028 13126
rect 5184 12434 5212 14826
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5276 13394 5304 13874
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5368 13258 5396 13806
rect 5644 13326 5672 14962
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5736 14385 5764 14894
rect 5722 14376 5778 14385
rect 5722 14311 5778 14320
rect 5920 14074 5948 14894
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5920 13870 5948 14010
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5632 13320 5684 13326
rect 5552 13268 5632 13274
rect 5552 13262 5684 13268
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5552 13246 5672 13262
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5000 12406 5120 12434
rect 5184 12406 5304 12434
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11898 5028 12038
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9897 4108 9998
rect 4436 9920 4488 9926
rect 4066 9888 4122 9897
rect 4436 9862 4488 9868
rect 4066 9823 4122 9832
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 9178 4016 9454
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 4080 8673 4108 9590
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4066 8664 4122 8673
rect 4066 8599 4122 8608
rect 3884 8560 3936 8566
rect 4172 8537 4200 9454
rect 4448 8974 4476 9862
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 3884 8502 3936 8508
rect 4158 8528 4214 8537
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3896 6905 3924 8502
rect 4158 8463 4214 8472
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5846 3280 6054
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3252 5642 3280 5782
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3160 5494 3280 5522
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4758 3188 5102
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3252 4570 3280 5494
rect 3160 4542 3280 4570
rect 3160 2990 3188 4542
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4146 3280 4422
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 3534 3280 3946
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3068 2746 3188 2774
rect 2962 2544 3018 2553
rect 2962 2479 3018 2488
rect 3160 800 3188 2746
rect 3252 2145 3280 2994
rect 3344 2774 3372 6258
rect 3988 6202 4016 7686
rect 4080 6866 4108 8298
rect 4264 8090 4292 8434
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4250 7712 4306 7721
rect 4250 7647 4306 7656
rect 4264 7546 4292 7647
rect 4356 7546 4384 8366
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6322 4108 6598
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3988 6174 4108 6202
rect 4080 6118 4108 6174
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3790 5808 3846 5817
rect 3790 5743 3846 5752
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 5370 3556 5646
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3436 4282 3464 5238
rect 3620 5166 3648 5510
rect 3804 5166 3832 5743
rect 4080 5710 4108 6054
rect 4172 5953 4200 6870
rect 4158 5944 4214 5953
rect 4158 5879 4214 5888
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3988 5030 4016 5646
rect 4080 5370 4108 5646
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4264 5234 4292 7346
rect 4342 6216 4398 6225
rect 4342 6151 4398 6160
rect 4252 5228 4304 5234
rect 4172 5188 4252 5216
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3606 4720 3662 4729
rect 3606 4655 3662 4664
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3620 4010 3648 4655
rect 3974 4176 4030 4185
rect 3884 4140 3936 4146
rect 4172 4146 4200 5188
rect 4252 5170 4304 5176
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 4282 4292 4422
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4356 4214 4384 6151
rect 4448 4622 4476 8774
rect 4540 8566 4568 9318
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6322 4568 6598
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4526 6080 4582 6089
rect 4526 6015 4582 6024
rect 4540 5778 4568 6015
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4632 4826 4660 11698
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 9994 4844 11018
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10810 4936 10950
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5000 9761 5028 9862
rect 4986 9752 5042 9761
rect 4986 9687 5042 9696
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 9489 5028 9522
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4724 9042 4752 9318
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 5234 4752 7822
rect 4908 7546 4936 8230
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5000 7478 5028 9318
rect 4988 7472 5040 7478
rect 4802 7440 4858 7449
rect 4988 7414 5040 7420
rect 4802 7375 4858 7384
rect 4816 7342 4844 7375
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5000 7002 5028 7278
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4908 6202 4936 6870
rect 4908 6174 5028 6202
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5370 4844 5510
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4436 4616 4488 4622
rect 4488 4576 4660 4604
rect 4436 4558 4488 4564
rect 4434 4312 4490 4321
rect 4434 4247 4490 4256
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 3974 4111 4030 4120
rect 4160 4140 4212 4146
rect 3884 4082 3936 4088
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3436 3534 3464 3878
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3698 3496 3754 3505
rect 3698 3431 3754 3440
rect 3422 3088 3478 3097
rect 3712 3058 3740 3431
rect 3422 3023 3478 3032
rect 3700 3052 3752 3058
rect 3436 2990 3464 3023
rect 3700 2994 3752 3000
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3344 2746 3464 2774
rect 3238 2136 3294 2145
rect 3238 2071 3294 2080
rect 3436 1442 3464 2746
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3436 1414 3556 1442
rect 3528 800 3556 1414
rect 3896 800 3924 4082
rect 3988 4010 4016 4111
rect 4160 4082 4212 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 3988 2514 4016 2751
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4080 2378 4108 4014
rect 4264 3913 4292 4082
rect 4448 4010 4476 4247
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4250 3904 4306 3913
rect 4250 3839 4306 3848
rect 4342 3496 4398 3505
rect 4342 3431 4398 3440
rect 4356 2446 4384 3431
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4080 1737 4108 1838
rect 4066 1728 4122 1737
rect 4066 1663 4122 1672
rect 4264 800 4292 2314
rect 4632 800 4660 4576
rect 4816 4128 4844 5170
rect 4724 4100 4844 4128
rect 4724 3890 4752 4100
rect 4802 4040 4858 4049
rect 4802 3975 4804 3984
rect 4856 3975 4858 3984
rect 4804 3946 4856 3952
rect 4724 3862 4844 3890
rect 4710 3768 4766 3777
rect 4710 3703 4712 3712
rect 4764 3703 4766 3712
rect 4712 3674 4764 3680
rect 4816 2582 4844 3862
rect 4908 3534 4936 6054
rect 5000 5030 5028 6174
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5092 4486 5120 12406
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5184 9518 5212 10066
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5184 8498 5212 9454
rect 5276 9450 5304 12406
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11830 5396 12038
rect 5460 11898 5488 13126
rect 5552 12102 5580 13246
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5644 11694 5672 12650
rect 5736 12442 5764 12718
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11762 5948 12038
rect 6012 11898 6040 15370
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6288 13394 6316 13942
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6564 12442 6592 16526
rect 6840 16454 6868 17614
rect 7300 17338 7328 19314
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6932 15162 6960 16458
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6840 12918 6868 13330
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5632 11688 5684 11694
rect 5630 11656 5632 11665
rect 5684 11656 5686 11665
rect 5630 11591 5686 11600
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8634 5304 8774
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5184 7274 5212 7890
rect 5276 7546 5304 7890
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 5794 5212 6598
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5914 5304 6190
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5184 5766 5304 5794
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5078 4312 5134 4321
rect 5078 4247 5134 4256
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4816 1902 4844 2382
rect 4804 1896 4856 1902
rect 4804 1838 4856 1844
rect 5000 800 5028 4150
rect 5092 4146 5120 4247
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5184 4010 5212 5510
rect 5276 5370 5304 5766
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5368 5250 5396 10406
rect 5460 8072 5488 10542
rect 5736 10062 5764 10610
rect 5828 10198 5856 11154
rect 6564 11121 6592 12038
rect 6656 11898 6684 12718
rect 6932 12714 6960 13126
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6932 12238 6960 12650
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6550 11112 6606 11121
rect 6550 11047 6606 11056
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6012 10266 6040 10950
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5552 9586 5580 9930
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 8673 5672 8774
rect 5630 8664 5686 8673
rect 5630 8599 5686 8608
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5460 8044 5580 8072
rect 5552 7954 5580 8044
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 7721 5580 7890
rect 5538 7712 5594 7721
rect 5538 7647 5594 7656
rect 5446 7576 5502 7585
rect 5446 7511 5502 7520
rect 5540 7540 5592 7546
rect 5460 7478 5488 7511
rect 5540 7482 5592 7488
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5276 5222 5396 5250
rect 5276 5098 5304 5222
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5368 5001 5396 5102
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5078 3496 5134 3505
rect 5078 3431 5134 3440
rect 5092 3194 5120 3431
rect 5276 3398 5304 4558
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5368 800 5396 4490
rect 5460 4049 5488 7142
rect 5552 6769 5580 7482
rect 5644 6934 5672 8366
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5538 6760 5594 6769
rect 5736 6746 5764 8298
rect 5538 6695 5594 6704
rect 5644 6718 5764 6746
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5552 6118 5580 6394
rect 5644 6338 5672 6718
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6458 5764 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5644 6310 5764 6338
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 4622 5580 5510
rect 5644 5234 5672 6122
rect 5736 5574 5764 6310
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5644 4214 5672 4966
rect 5828 4570 5856 8298
rect 5920 7177 5948 9862
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6564 9625 6592 10950
rect 6656 10742 6684 11154
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6734 10840 6790 10849
rect 6734 10775 6790 10784
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6748 10577 6776 10775
rect 6932 10674 6960 10950
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6734 10568 6790 10577
rect 6734 10503 6790 10512
rect 6918 10568 6974 10577
rect 6918 10503 6920 10512
rect 6972 10503 6974 10512
rect 6920 10474 6972 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6550 9616 6606 9625
rect 6550 9551 6606 9560
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5906 7168 5962 7177
rect 5906 7103 5962 7112
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 6254 5948 6666
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5920 5166 5948 5306
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4729 5948 4966
rect 5906 4720 5962 4729
rect 5906 4655 5962 4664
rect 5736 4542 5856 4570
rect 5736 4321 5764 4542
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5722 4312 5778 4321
rect 5722 4247 5778 4256
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5446 4040 5502 4049
rect 5446 3975 5502 3984
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5552 3738 5580 3946
rect 5630 3904 5686 3913
rect 5630 3839 5686 3848
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 2038 5488 3402
rect 5538 3224 5594 3233
rect 5538 3159 5540 3168
rect 5592 3159 5594 3168
rect 5540 3130 5592 3136
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5552 2106 5580 2382
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 5644 1442 5672 3839
rect 5736 1562 5764 4247
rect 5828 3738 5856 4422
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5920 3913 5948 4014
rect 5906 3904 5962 3913
rect 5906 3839 5962 3848
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 6012 3618 6040 8842
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6380 6798 6408 7346
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6460 6452 6512 6458
rect 6656 6440 6684 9415
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 7041 6776 8842
rect 6840 8129 6868 10406
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9654 6960 9862
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6932 9178 6960 9454
rect 7024 9450 7052 14826
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 13410 7144 14350
rect 7208 13530 7236 16526
rect 7484 16454 7512 18226
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 15502 7696 15982
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7392 14074 7420 14894
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7116 13382 7236 13410
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7116 12238 7144 12718
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 11082 7144 11630
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7116 8401 7144 9930
rect 7102 8392 7158 8401
rect 6920 8356 6972 8362
rect 7102 8327 7158 8336
rect 6920 8298 6972 8304
rect 6826 8120 6882 8129
rect 6826 8055 6882 8064
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6734 7032 6790 7041
rect 6840 7002 6868 7754
rect 6734 6967 6790 6976
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6458 6776 6598
rect 6512 6412 6684 6440
rect 6736 6452 6788 6458
rect 6460 6394 6512 6400
rect 6736 6394 6788 6400
rect 6472 6186 6500 6394
rect 6460 6180 6512 6186
rect 6460 6122 6512 6128
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6564 5817 6592 6122
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6550 5808 6606 5817
rect 6460 5772 6512 5778
rect 6550 5743 6606 5752
rect 6460 5714 6512 5720
rect 6472 5658 6500 5714
rect 6472 5630 6592 5658
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6564 5370 6592 5630
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6104 4554 6132 5306
rect 6748 5216 6776 6054
rect 6840 5914 6868 6802
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6748 5188 6868 5216
rect 6734 5128 6790 5137
rect 6734 5063 6736 5072
rect 6788 5063 6790 5072
rect 6736 5034 6788 5040
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4690 6408 4966
rect 6748 4706 6776 5034
rect 6840 4826 6868 5188
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6564 4678 6776 4706
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 6090 3904 6146 3913
rect 6090 3839 6146 3848
rect 5828 3590 6040 3618
rect 6104 3602 6132 3839
rect 6092 3596 6144 3602
rect 5828 2446 5856 3590
rect 6092 3538 6144 3544
rect 6104 3466 6132 3538
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6196 3398 6224 4150
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6288 3738 6316 4082
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6288 3602 6316 3674
rect 6564 3602 6592 4678
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6656 3534 6684 4422
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5920 2774 5948 3334
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 5998 2952 6054 2961
rect 5998 2887 6000 2896
rect 6052 2887 6054 2896
rect 6000 2858 6052 2864
rect 5920 2746 6040 2774
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5828 1834 5856 2382
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 1873 5948 2246
rect 5906 1864 5962 1873
rect 5816 1828 5868 1834
rect 5906 1799 5962 1808
rect 5816 1770 5868 1776
rect 5724 1556 5776 1562
rect 5724 1498 5776 1504
rect 6012 1442 6040 2746
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 5644 1414 5764 1442
rect 6012 1414 6132 1442
rect 5736 800 5764 1414
rect 6104 800 6132 1414
rect 6472 800 6500 1498
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6564 762 6592 3402
rect 6748 2990 6776 4558
rect 6840 3738 6868 4762
rect 6932 4214 6960 8298
rect 7208 7546 7236 13382
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7300 10266 7328 12038
rect 7392 11898 7420 12038
rect 7484 11898 7512 15438
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8312 14074 8340 14282
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7852 12986 7880 13398
rect 8128 13326 8156 13942
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8116 13320 8168 13326
rect 8220 13297 8248 13330
rect 8116 13262 8168 13268
rect 8206 13288 8262 13297
rect 8206 13223 8262 13232
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7286 10024 7342 10033
rect 7286 9959 7342 9968
rect 7300 7886 7328 9959
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7576 9722 7604 9862
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7668 9586 7696 9862
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 8838 7604 9318
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7392 7478 7420 8774
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 6633 7052 7278
rect 7102 6896 7158 6905
rect 7102 6831 7158 6840
rect 7010 6624 7066 6633
rect 7010 6559 7066 6568
rect 7024 6186 7052 6559
rect 7116 6497 7144 6831
rect 7484 6794 7512 8230
rect 7576 8090 7604 8366
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7668 7290 7696 8978
rect 7760 8945 7788 12106
rect 7852 11558 7880 12922
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12442 8064 12718
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8036 12170 8064 12378
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 9908 7880 11494
rect 7944 11257 7972 12038
rect 7930 11248 7986 11257
rect 7930 11183 7986 11192
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 10130 8064 11154
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7932 9920 7984 9926
rect 7852 9880 7932 9908
rect 7932 9862 7984 9868
rect 8036 9625 8064 10066
rect 8022 9616 8078 9625
rect 8022 9551 8078 9560
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7746 8936 7802 8945
rect 7746 8871 7802 8880
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7576 7262 7696 7290
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7480 6788 7532 6794
rect 7208 6718 7420 6746
rect 7480 6730 7532 6736
rect 7102 6488 7158 6497
rect 7102 6423 7158 6432
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7116 5681 7144 6258
rect 7102 5672 7158 5681
rect 7102 5607 7158 5616
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3194 6960 4014
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6826 2680 6882 2689
rect 6826 2615 6882 2624
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6656 2281 6684 2518
rect 6840 2446 6868 2615
rect 7024 2446 7052 4966
rect 7208 4604 7236 6718
rect 7392 6662 7420 6718
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7116 4576 7236 4604
rect 7116 3482 7144 4576
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7208 4049 7236 4082
rect 7194 4040 7250 4049
rect 7194 3975 7250 3984
rect 7116 3454 7236 3482
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3058 7144 3334
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7208 2938 7236 3454
rect 7300 3126 7328 6598
rect 7576 6338 7604 7262
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7484 6310 7604 6338
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5545 7420 6190
rect 7378 5536 7434 5545
rect 7378 5471 7434 5480
rect 7392 5001 7420 5471
rect 7378 4992 7434 5001
rect 7378 4927 7434 4936
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 3194 7420 4422
rect 7484 4146 7512 6310
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 4282 7604 6122
rect 7668 4622 7696 7142
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7470 3632 7526 3641
rect 7470 3567 7526 3576
rect 7484 3534 7512 3567
rect 7576 3534 7604 4218
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7562 3224 7618 3233
rect 7380 3188 7432 3194
rect 7562 3159 7618 3168
rect 7380 3130 7432 3136
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7116 2910 7236 2938
rect 7576 2922 7604 3159
rect 7564 2916 7616 2922
rect 7116 2514 7144 2910
rect 7564 2858 7616 2864
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6828 2440 6880 2446
rect 6734 2408 6790 2417
rect 6828 2382 6880 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6734 2343 6790 2352
rect 6748 2310 6776 2343
rect 6736 2304 6788 2310
rect 6642 2272 6698 2281
rect 6736 2246 6788 2252
rect 6642 2207 6698 2216
rect 7116 1698 7144 2450
rect 7104 1692 7156 1698
rect 7104 1634 7156 1640
rect 6748 870 6868 898
rect 6748 762 6776 870
rect 6840 800 6868 870
rect 7208 800 7236 2790
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 1970 7512 2246
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7576 800 7604 2858
rect 7668 2854 7696 4082
rect 7760 2854 7788 7278
rect 7852 6905 7880 7890
rect 7838 6896 7894 6905
rect 7838 6831 7894 6840
rect 7944 5794 7972 9046
rect 8128 7818 8156 12242
rect 8220 12238 8248 12650
rect 8496 12442 8524 16526
rect 8588 16454 8616 19314
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9324 14618 9352 15302
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9416 14074 9444 17614
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9692 14278 9720 14554
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9784 13841 9812 14214
rect 10336 14074 10364 14214
rect 10428 14074 10456 19790
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 9770 13832 9826 13841
rect 8576 13796 8628 13802
rect 9770 13767 9826 13776
rect 10140 13796 10192 13802
rect 8576 13738 8628 13744
rect 10140 13738 10192 13744
rect 8588 13530 8616 13738
rect 10152 13705 10180 13738
rect 10138 13696 10194 13705
rect 8747 13628 9055 13637
rect 10138 13631 10194 13640
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 10230 13288 10286 13297
rect 10230 13223 10286 13232
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 9140 12102 9168 12786
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9586 12336 9642 12345
rect 9586 12271 9588 12280
rect 9640 12271 9642 12280
rect 9588 12242 9640 12248
rect 9692 12238 9720 12718
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11762 9168 12038
rect 9876 11898 9904 12106
rect 9968 11898 9996 12310
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9232 11801 9260 11834
rect 9218 11792 9274 11801
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9128 11756 9180 11762
rect 9218 11727 9274 11736
rect 9128 11698 9180 11704
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8220 11014 8248 11222
rect 8680 11218 8708 11698
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 9140 11150 9168 11698
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8944 10736 8996 10742
rect 8942 10704 8944 10713
rect 8996 10704 8998 10713
rect 8942 10639 8998 10648
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 10033 8248 10066
rect 8206 10024 8262 10033
rect 8206 9959 8262 9968
rect 8312 8514 8340 10406
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9654 8432 9862
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8634 8432 8774
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8312 8486 8432 8514
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 8022 8340 8366
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7546 8248 7686
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8036 5817 8064 7414
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 7041 8248 7142
rect 8206 7032 8262 7041
rect 8312 7002 8340 7346
rect 8206 6967 8262 6976
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7852 5766 7972 5794
rect 8022 5808 8078 5817
rect 7852 5710 7880 5766
rect 8022 5743 8078 5752
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7944 5302 7972 5578
rect 8128 5370 8156 6394
rect 8220 6225 8248 6802
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8206 6216 8262 6225
rect 8206 6151 8262 6160
rect 8312 5930 8340 6598
rect 8220 5902 8340 5930
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7840 4480 7892 4486
rect 8128 4457 8156 4966
rect 7840 4422 7892 4428
rect 8114 4448 8170 4457
rect 7852 4185 7880 4422
rect 8114 4383 8170 4392
rect 7838 4176 7894 4185
rect 7838 4111 7894 4120
rect 8220 4026 8248 5902
rect 8300 5840 8352 5846
rect 8298 5808 8300 5817
rect 8352 5808 8354 5817
rect 8298 5743 8354 5752
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5409 8340 5510
rect 8298 5400 8354 5409
rect 8298 5335 8354 5344
rect 8404 4842 8432 8486
rect 8496 5234 8524 8570
rect 8680 8498 8708 8910
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 8424 8628 8430
rect 8772 8378 8800 8774
rect 8576 8366 8628 8372
rect 8588 8090 8616 8366
rect 8680 8350 8800 8378
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8680 6474 8708 8350
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7585 8984 7686
rect 8942 7576 8998 7585
rect 8942 7511 8998 7520
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8588 6446 8708 6474
rect 9048 6458 9076 6598
rect 9036 6452 9088 6458
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8588 5114 8616 6446
rect 9036 6394 9088 6400
rect 8668 6384 8720 6390
rect 8666 6352 8668 6361
rect 8720 6352 8722 6361
rect 8666 6287 8722 6296
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8760 5908 8812 5914
rect 8812 5868 9076 5896
rect 8760 5850 8812 5856
rect 9048 5778 9076 5868
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9140 5166 9168 9318
rect 9324 6390 9352 10610
rect 10244 10470 10272 13223
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9761 9444 9862
rect 9402 9752 9458 9761
rect 9402 9687 9458 9696
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8634 9536 8774
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9692 7478 9720 10066
rect 9876 9654 9904 10406
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 9722 9996 9862
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9784 7886 9812 9007
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9876 8090 9904 8366
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9416 6798 9444 7278
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9956 6656 10008 6662
rect 9954 6624 9956 6633
rect 10008 6624 10010 6633
rect 9954 6559 10010 6568
rect 9968 6390 9996 6559
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 10152 6202 10180 7278
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 6322 10272 7142
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9324 5710 9352 6190
rect 10152 6174 10272 6202
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 9508 5914 9536 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9678 5536 9734 5545
rect 9678 5471 9734 5480
rect 8496 5086 8616 5114
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 8496 5001 8524 5086
rect 8576 5024 8628 5030
rect 8482 4992 8538 5001
rect 8576 4966 8628 4972
rect 8482 4927 8538 4936
rect 8404 4814 8524 4842
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8128 3998 8248 4026
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7852 3074 7880 3538
rect 7852 3046 7972 3074
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7668 1494 7696 2246
rect 7852 1766 7880 2926
rect 7944 2446 7972 3046
rect 8036 2922 8064 3878
rect 8128 3602 8156 3998
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 8128 3194 8156 3431
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8114 3088 8170 3097
rect 8114 3023 8170 3032
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 8128 2650 8156 3023
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7944 2310 7972 2382
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 8220 1766 8248 3878
rect 8312 3738 8340 4558
rect 8404 4185 8432 4626
rect 8390 4176 8446 4185
rect 8390 4111 8446 4120
rect 8496 4026 8524 4814
rect 8404 3998 8524 4026
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8298 3632 8354 3641
rect 8298 3567 8354 3576
rect 8312 2106 8340 3567
rect 8404 3058 8432 3998
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8496 2514 8524 3878
rect 8588 3534 8616 4966
rect 8680 3720 8708 5102
rect 9692 5030 9720 5471
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 9218 4448 9274 4457
rect 8864 4078 8892 4422
rect 9218 4383 9274 4392
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8852 3732 8904 3738
rect 8680 3692 8800 3720
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8680 3369 8708 3538
rect 8666 3360 8722 3369
rect 8666 3295 8722 3304
rect 8668 2984 8720 2990
rect 8772 2972 8800 3692
rect 8852 3674 8904 3680
rect 8864 3194 8892 3674
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8956 3126 8984 3606
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9048 3369 9076 3470
rect 9034 3360 9090 3369
rect 9034 3295 9090 3304
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8720 2944 8800 2972
rect 8668 2926 8720 2932
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8300 2100 8352 2106
rect 9140 2088 9168 4082
rect 9232 3058 9260 4383
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9324 3641 9352 3946
rect 9310 3632 9366 3641
rect 9416 3602 9444 4966
rect 9494 4584 9550 4593
rect 9494 4519 9550 4528
rect 9508 4486 9536 4519
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9494 4312 9550 4321
rect 9494 4247 9550 4256
rect 9508 3777 9536 4247
rect 9692 4214 9720 4422
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9784 4146 9812 6054
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9770 4040 9826 4049
rect 9770 3975 9826 3984
rect 9494 3768 9550 3777
rect 9494 3703 9550 3712
rect 9784 3670 9812 3975
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9310 3567 9366 3576
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3504 9640 3510
rect 9588 3446 9640 3452
rect 9496 3392 9548 3398
rect 9310 3360 9366 3369
rect 9310 3295 9366 3304
rect 9416 3352 9496 3380
rect 9324 3194 9352 3295
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9232 2802 9260 2858
rect 9416 2802 9444 3352
rect 9496 3334 9548 3340
rect 9494 3224 9550 3233
rect 9494 3159 9496 3168
rect 9548 3159 9550 3168
rect 9496 3130 9548 3136
rect 9232 2774 9444 2802
rect 9218 2680 9274 2689
rect 9218 2615 9274 2624
rect 9232 2582 9260 2615
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9600 2446 9628 3446
rect 9692 3058 9720 3538
rect 9784 3233 9812 3606
rect 9770 3224 9826 3233
rect 9770 3159 9826 3168
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9678 2544 9734 2553
rect 9678 2479 9734 2488
rect 9692 2446 9720 2479
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 8300 2042 8352 2048
rect 9048 2060 9168 2088
rect 7840 1760 7892 1766
rect 7840 1702 7892 1708
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 7932 1692 7984 1698
rect 7932 1634 7984 1640
rect 7656 1488 7708 1494
rect 7656 1430 7708 1436
rect 7944 800 7972 1634
rect 8312 800 8340 2042
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 8680 800 8708 1770
rect 9048 800 9076 2060
rect 9416 800 9444 2246
rect 9692 1426 9720 2246
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9784 800 9812 2926
rect 9876 2582 9904 5850
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5370 9996 5510
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9956 5024 10008 5030
rect 9954 4992 9956 5001
rect 10008 4992 10010 5001
rect 9954 4927 10010 4936
rect 9954 4040 10010 4049
rect 9954 3975 9956 3984
rect 10008 3975 10010 3984
rect 9956 3946 10008 3952
rect 10060 2774 10088 5170
rect 10152 3097 10180 6054
rect 10244 3534 10272 6174
rect 10336 4622 10364 7686
rect 10428 7290 10456 12718
rect 10520 8974 10548 14350
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 14074 10824 14214
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11286 10640 12038
rect 10600 11280 10652 11286
rect 10704 11257 10732 13126
rect 10888 12434 10916 14418
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 10968 13864 11020 13870
rect 11152 13864 11204 13870
rect 11020 13812 11152 13818
rect 10968 13806 11204 13812
rect 10980 13790 11192 13806
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11072 12986 11100 13398
rect 11716 13394 11744 14554
rect 11978 13968 12034 13977
rect 11888 13932 11940 13938
rect 11978 13903 11980 13912
rect 11888 13874 11940 13880
rect 12032 13903 12034 13912
rect 11980 13874 12032 13880
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 13258 11744 13330
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11808 12442 11836 13466
rect 11900 13462 11928 13874
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11796 12436 11848 12442
rect 10888 12406 11008 12434
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11222 10652 11228
rect 10690 11248 10746 11257
rect 10612 9586 10640 11222
rect 10690 11183 10746 11192
rect 10692 11144 10744 11150
rect 10796 11121 10824 12038
rect 10980 11150 11008 12406
rect 11796 12378 11848 12384
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10968 11144 11020 11150
rect 10692 11086 10744 11092
rect 10782 11112 10838 11121
rect 10704 10062 10732 11086
rect 10968 11086 11020 11092
rect 10782 11047 10838 11056
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 11072 9722 11100 12242
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11716 11762 11744 12174
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11164 9994 11192 10746
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10428 7262 10548 7290
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10138 3088 10194 3097
rect 10138 3023 10194 3032
rect 9968 2746 10088 2774
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 6564 734 6776 762
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 9876 762 9904 2518
rect 9968 1426 9996 2746
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10060 2038 10088 2246
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 10428 1902 10456 7142
rect 10520 3942 10548 7262
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10612 3058 10640 8774
rect 10888 8401 10916 9454
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10874 8392 10930 8401
rect 10874 8327 10930 8336
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7546 10732 7686
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10980 6662 11008 8502
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10690 6488 10746 6497
rect 10690 6423 10746 6432
rect 10704 4146 10732 6423
rect 10782 6216 10838 6225
rect 10782 6151 10838 6160
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 3534 10732 4082
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10796 3466 10824 6151
rect 10980 5574 11008 6598
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10876 4616 10928 4622
rect 10980 4593 11008 4626
rect 10876 4558 10928 4564
rect 10966 4584 11022 4593
rect 10888 4146 10916 4558
rect 11072 4554 11100 9454
rect 11256 9382 11284 11698
rect 11794 11384 11850 11393
rect 11794 11319 11850 11328
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11336 9172 11388 9178
rect 11256 9132 11336 9160
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8634 11192 8910
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 6866 11192 8570
rect 11256 7954 11284 9132
rect 11336 9114 11388 9120
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11716 8242 11744 9930
rect 11808 9178 11836 11319
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8362 11836 8774
rect 11900 8566 11928 10202
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11888 8424 11940 8430
rect 11886 8392 11888 8401
rect 11940 8392 11942 8401
rect 11796 8356 11848 8362
rect 11886 8327 11942 8336
rect 11796 8298 11848 8304
rect 11716 8214 11928 8242
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11242 7848 11298 7857
rect 11242 7783 11298 7792
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11164 6458 11192 6802
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11164 5914 11192 6394
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11164 5234 11192 5850
rect 11256 5681 11284 7783
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11716 7546 11744 7890
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11716 6458 11744 6734
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4690 11192 5170
rect 11716 5166 11744 6258
rect 11900 6118 11928 8214
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 10966 4519 11022 4528
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10416 1896 10468 1902
rect 10416 1838 10468 1844
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 10060 870 10180 898
rect 10060 762 10088 870
rect 10152 800 10180 870
rect 10520 800 10548 2994
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 10704 1902 10732 2246
rect 10692 1896 10744 1902
rect 10692 1838 10744 1844
rect 10888 800 10916 4082
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 2145 11008 2246
rect 10966 2136 11022 2145
rect 10966 2071 11022 2080
rect 11072 1306 11100 3946
rect 11164 3602 11192 4626
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 3058 11192 3538
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 2650 11192 2994
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2582 11284 4490
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11532 4010 11560 4082
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3670 11376 3878
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11716 2446 11744 4966
rect 11808 2514 11836 6054
rect 11886 5536 11942 5545
rect 11886 5471 11942 5480
rect 11900 5370 11928 5471
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11886 5264 11942 5273
rect 11886 5199 11942 5208
rect 11900 4049 11928 5199
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11900 3942 11928 3975
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11992 2774 12020 13738
rect 12084 13530 12112 16662
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12176 12986 12204 17138
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 20732 16658 20760 17478
rect 21284 17241 21312 17478
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12084 8906 12112 12854
rect 12268 12434 12296 15506
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 14074 12940 14214
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12176 12406 12296 12434
rect 12176 12102 12204 12406
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12176 11354 12204 12038
rect 12268 11558 12296 12106
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 9586 12204 11018
rect 12268 10674 12296 11494
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10062 12296 10610
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12268 9926 12296 9998
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12254 9616 12310 9625
rect 12164 9580 12216 9586
rect 12254 9551 12310 9560
rect 12164 9522 12216 9528
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12084 8362 12112 8842
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7750 12204 8230
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12268 7528 12296 9551
rect 12176 7500 12296 7528
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 5352 12112 7346
rect 12176 6322 12204 7500
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12084 5324 12204 5352
rect 12070 5264 12126 5273
rect 12070 5199 12126 5208
rect 12084 5001 12112 5199
rect 12070 4992 12126 5001
rect 12070 4927 12126 4936
rect 12176 4842 12204 5324
rect 12084 4814 12204 4842
rect 12084 3913 12112 4814
rect 12360 4672 12388 13806
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12440 9648 12492 9654
rect 12438 9616 12440 9625
rect 12492 9616 12494 9625
rect 12438 9551 12494 9560
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12452 5250 12480 7482
rect 12544 5386 12572 13126
rect 13004 12434 13032 13670
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12986 13124 13126
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13176 12436 13228 12442
rect 13004 12406 13124 12434
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12728 10713 12756 11222
rect 12714 10704 12770 10713
rect 12714 10639 12770 10648
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 7818 12664 9318
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12624 7404 12676 7410
rect 12728 7392 12756 10639
rect 13096 10470 13124 12406
rect 13176 12378 13228 12384
rect 13188 12102 13216 12378
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13188 11150 13216 11698
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13004 10198 13032 10406
rect 12992 10192 13044 10198
rect 13280 10146 13308 14554
rect 13818 13696 13874 13705
rect 13818 13631 13874 13640
rect 13832 12442 13860 13631
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13372 11082 13400 11766
rect 14292 11762 14320 12038
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 13464 11558 13492 11591
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13740 11218 13768 11698
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 12992 10134 13044 10140
rect 13188 10118 13308 10146
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9568 12848 9862
rect 12900 9580 12952 9586
rect 12820 9540 12900 9568
rect 12820 8974 12848 9540
rect 12900 9522 12952 9528
rect 13188 9450 13216 10118
rect 13266 10024 13322 10033
rect 13266 9959 13322 9968
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12820 8514 12848 8910
rect 12992 8900 13044 8906
rect 13044 8860 13124 8888
rect 12992 8842 13044 8848
rect 12820 8498 13032 8514
rect 12820 8492 13044 8498
rect 12820 8486 12992 8492
rect 12820 7886 12848 8486
rect 12992 8434 13044 8440
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7410 12848 7822
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12676 7364 12756 7392
rect 12808 7404 12860 7410
rect 12624 7346 12676 7352
rect 12808 7346 12860 7352
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12544 5358 12756 5386
rect 12452 5234 12664 5250
rect 12452 5228 12676 5234
rect 12452 5222 12624 5228
rect 12624 5170 12676 5176
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12176 4644 12388 4672
rect 12176 4282 12204 4644
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12360 4282 12388 4490
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4282 12480 4422
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12070 3904 12126 3913
rect 12070 3839 12126 3848
rect 12544 3466 12572 4694
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 11992 2746 12112 2774
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11612 1624 11664 1630
rect 11612 1566 11664 1572
rect 11072 1278 11284 1306
rect 11256 800 11284 1278
rect 11624 800 11652 1566
rect 9876 734 10088 762
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11716 762 11744 2382
rect 11808 1630 11836 2450
rect 12084 1873 12112 2746
rect 12070 1864 12126 1873
rect 12070 1799 12126 1808
rect 12072 1760 12124 1766
rect 12072 1702 12124 1708
rect 11796 1624 11848 1630
rect 11796 1566 11848 1572
rect 12084 1494 12112 1702
rect 12072 1488 12124 1494
rect 12072 1430 12124 1436
rect 11900 870 12020 898
rect 11900 762 11928 870
rect 11992 800 12020 870
rect 12360 800 12388 3130
rect 12728 2774 12756 5358
rect 12820 4622 12848 6326
rect 12912 4826 12940 7754
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 13096 4162 13124 8860
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13188 7274 13216 8502
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13188 6934 13216 7210
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13188 6322 13216 6394
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 12820 4134 13124 4162
rect 13280 4146 13308 9959
rect 13372 8634 13400 11018
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 8634 13492 10406
rect 13832 8974 13860 11494
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 14278 8936 14334 8945
rect 14278 8871 14334 8880
rect 14292 8838 14320 8871
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13726 8528 13782 8537
rect 13726 8463 13728 8472
rect 13780 8463 13782 8472
rect 13728 8434 13780 8440
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13372 5914 13400 6258
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13648 5914 13676 6190
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13372 5778 13400 5850
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13372 5370 13400 5714
rect 13740 5710 13768 6054
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13832 5574 13860 6054
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14292 5642 14320 8774
rect 14384 7818 14412 12106
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9654 14780 10406
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14660 6662 14688 8842
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15212 8498 15240 8570
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15304 7546 15332 8366
rect 15396 8090 15424 15030
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15580 11898 15608 14894
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 15672 12102 15700 13670
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16776 12170 16804 12718
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15488 10674 15516 11290
rect 15580 11150 15608 11834
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15672 10810 15700 12038
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16500 11354 16528 11630
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15580 9042 15608 9590
rect 15750 9480 15806 9489
rect 15750 9415 15806 9424
rect 15764 9382 15792 9415
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15580 8634 15608 8978
rect 15764 8838 15792 9318
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15856 8294 15884 10610
rect 16304 10600 16356 10606
rect 15934 10568 15990 10577
rect 16304 10542 16356 10548
rect 15934 10503 15990 10512
rect 15948 9178 15976 10503
rect 16316 9926 16344 10542
rect 16408 10470 16436 11018
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16670 10160 16726 10169
rect 16670 10095 16726 10104
rect 16684 9994 16712 10095
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9654 16344 9862
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 17052 9450 17080 11018
rect 17328 10266 17356 12106
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17788 10577 17816 10610
rect 17774 10568 17830 10577
rect 17774 10503 17830 10512
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 17880 8634 17908 13330
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11830 18368 12038
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 9625 18184 11494
rect 18248 10810 18276 11698
rect 18340 11694 18368 11766
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18340 11150 18368 11630
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18432 10062 18460 12582
rect 18984 11898 19012 13670
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19064 12436 19116 12442
rect 19720 12434 19748 13262
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12646 20760 13126
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 19720 12406 19840 12434
rect 19064 12378 19116 12384
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18984 11082 19012 11834
rect 19076 11354 19104 12378
rect 19812 11558 19840 12406
rect 20536 12232 20588 12238
rect 20534 12200 20536 12209
rect 20588 12200 20590 12209
rect 20732 12170 20760 12582
rect 20810 12336 20866 12345
rect 20810 12271 20866 12280
rect 20534 12135 20590 12144
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20824 11830 20852 12271
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 19800 11552 19852 11558
rect 20824 11506 20852 11766
rect 19800 11494 19852 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 19812 10674 19840 11494
rect 20732 11478 20852 11506
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19076 10266 19104 10406
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19260 9654 19288 9930
rect 19352 9722 19380 9930
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 9648 19300 9654
rect 18142 9616 18198 9625
rect 19248 9590 19300 9596
rect 18142 9551 18144 9560
rect 18196 9551 18198 9560
rect 18420 9580 18472 9586
rect 18144 9522 18196 9528
rect 18420 9522 18472 9528
rect 18156 9491 18184 9522
rect 18432 9178 18460 9522
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15856 7750 15884 7958
rect 15948 7954 15976 8570
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17314 8392 17370 8401
rect 17314 8327 17370 8336
rect 17328 8090 17356 8327
rect 17604 8090 17632 8502
rect 17316 8084 17368 8090
rect 17592 8084 17644 8090
rect 17368 8044 17448 8072
rect 17316 8026 17368 8032
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15948 7546 15976 7890
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 7002 16252 7210
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15750 6760 15806 6769
rect 15200 6724 15252 6730
rect 15750 6695 15752 6704
rect 15200 6666 15252 6672
rect 15804 6695 15806 6704
rect 15752 6666 15804 6672
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6338 14688 6598
rect 14660 6322 14872 6338
rect 15212 6322 15240 6666
rect 14660 6316 14884 6322
rect 14660 6310 14832 6316
rect 14832 6258 14884 6264
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 15566 5808 15622 5817
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14384 5574 14412 5782
rect 14464 5772 14516 5778
rect 15566 5743 15622 5752
rect 14464 5714 14516 5720
rect 13820 5568 13872 5574
rect 14096 5568 14148 5574
rect 13820 5510 13872 5516
rect 14094 5536 14096 5545
rect 14372 5568 14424 5574
rect 14148 5536 14150 5545
rect 14372 5510 14424 5516
rect 14094 5471 14150 5480
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 5234 13400 5306
rect 14108 5234 14136 5471
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13372 4826 13400 5170
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13726 4856 13782 4865
rect 13945 4859 14253 4868
rect 13360 4820 13412 4826
rect 13726 4791 13782 4800
rect 14280 4820 14332 4826
rect 13360 4762 13412 4768
rect 13372 4554 13400 4762
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13372 4214 13400 4490
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13268 4140 13320 4146
rect 12820 4010 12848 4134
rect 13268 4082 13320 4088
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12452 2746 12756 2774
rect 12452 1902 12480 2746
rect 12820 2446 12848 3946
rect 12912 3126 12940 4014
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13280 2922 13308 4082
rect 13556 3534 13584 4422
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13740 3058 13768 4791
rect 14280 4762 14332 4768
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14292 3670 14320 4762
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14280 3664 14332 3670
rect 14278 3632 14280 3641
rect 14332 3632 14334 3641
rect 14278 3567 14334 3576
rect 14384 3505 14412 4422
rect 14476 4214 14504 5714
rect 15580 5642 15608 5743
rect 15764 5642 15792 6666
rect 16040 6458 16068 6802
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16040 5914 16068 6394
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16040 5778 16068 5850
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15842 5672 15898 5681
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15752 5636 15804 5642
rect 15842 5607 15898 5616
rect 15752 5578 15804 5584
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14568 4593 14596 4966
rect 14554 4584 14610 4593
rect 14554 4519 14610 4528
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14568 3516 14596 4519
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 14648 3528 14700 3534
rect 14370 3496 14426 3505
rect 14568 3488 14648 3516
rect 14648 3470 14700 3476
rect 14370 3431 14426 3440
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13360 2984 13412 2990
rect 13358 2952 13360 2961
rect 13412 2952 13414 2961
rect 13268 2916 13320 2922
rect 13358 2887 13414 2896
rect 13268 2858 13320 2864
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12808 2304 12860 2310
rect 12728 2264 12808 2292
rect 12440 1896 12492 1902
rect 12440 1838 12492 1844
rect 12728 800 12756 2264
rect 12808 2246 12860 2252
rect 13096 800 13124 2518
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13188 2106 13216 2382
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13464 800 13492 2790
rect 13832 2514 13860 3334
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 800 13860 2314
rect 14108 1834 14136 2382
rect 14096 1828 14148 1834
rect 14096 1770 14148 1776
rect 14292 1442 14320 2790
rect 14384 2310 14412 2926
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14200 1414 14320 1442
rect 14200 800 14228 1414
rect 14568 800 14596 2518
rect 15028 2378 15056 3402
rect 15120 2514 15148 4218
rect 15580 3670 15608 5578
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15764 4554 15792 4966
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15856 3534 15884 5607
rect 16040 5370 16068 5714
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16040 4622 16068 5306
rect 16316 4758 16344 7754
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16408 7002 16436 7482
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16776 6662 16804 7142
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16960 5273 16988 6258
rect 17132 5296 17184 5302
rect 16946 5264 17002 5273
rect 17132 5238 17184 5244
rect 16946 5199 17002 5208
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16040 4214 16068 4558
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16028 4208 16080 4214
rect 16028 4150 16080 4156
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 3738 15976 4082
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16040 3602 16068 4150
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16408 3534 16436 3878
rect 16868 3738 16896 4218
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14936 800 14964 2246
rect 15212 2009 15240 2382
rect 15198 2000 15254 2009
rect 15198 1935 15254 1944
rect 15304 800 15332 2790
rect 15396 1766 15424 2994
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15384 1760 15436 1766
rect 15384 1702 15436 1708
rect 15672 800 15700 2790
rect 15844 2440 15896 2446
rect 15948 2417 15976 2994
rect 16408 2774 16436 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16856 3188 16908 3194
rect 16960 3176 16988 4626
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17052 3194 17080 4422
rect 17144 4049 17172 5238
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17130 4040 17186 4049
rect 17130 3975 17186 3984
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16908 3148 16988 3176
rect 17040 3188 17092 3194
rect 16856 3130 16908 3136
rect 17040 3130 17092 3136
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16408 2746 16620 2774
rect 16592 2650 16620 2746
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 15844 2382 15896 2388
rect 15934 2408 15990 2417
rect 15856 1970 15884 2382
rect 15934 2343 15990 2352
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 15844 1964 15896 1970
rect 15844 1906 15896 1912
rect 16040 800 16068 2246
rect 16408 800 16436 2518
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 1442 16988 2790
rect 17052 2038 17080 2926
rect 17040 2032 17092 2038
rect 17040 1974 17092 1980
rect 16776 1414 16988 1442
rect 16776 800 16804 1414
rect 17144 800 17172 3606
rect 17236 3097 17264 4082
rect 17328 3942 17356 6598
rect 17420 6322 17448 8044
rect 17592 8026 17644 8032
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17696 7546 17724 8026
rect 17972 7546 18000 8842
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18432 7886 18460 8434
rect 19536 8362 19564 9318
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 18512 8016 18564 8022
rect 18510 7984 18512 7993
rect 18564 7984 18566 7993
rect 18510 7919 18566 7928
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17696 7410 17724 7482
rect 17972 7449 18000 7482
rect 17958 7440 18014 7449
rect 17684 7404 17736 7410
rect 17958 7375 18014 7384
rect 17684 7346 17736 7352
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 5710 17632 6054
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 4282 17908 4422
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 17972 4010 18000 5578
rect 18064 5166 18092 6666
rect 18156 6458 18184 6802
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18142 5128 18198 5137
rect 18064 4185 18092 5102
rect 18142 5063 18198 5072
rect 18156 5030 18184 5063
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18050 4176 18106 4185
rect 18050 4111 18106 4120
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17222 3088 17278 3097
rect 17222 3023 17278 3032
rect 17512 800 17540 3334
rect 17788 2990 17816 3878
rect 18156 3754 18184 4966
rect 18248 4826 18276 5510
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 17972 3726 18184 3754
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 17880 800 17908 3130
rect 17972 2774 18000 3726
rect 18248 3618 18276 4762
rect 18156 3590 18276 3618
rect 18156 3466 18184 3590
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18248 2774 18276 3402
rect 18340 3126 18368 6598
rect 18524 5234 18552 7919
rect 19536 7478 19564 8298
rect 19628 8090 19656 10610
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19720 9178 19748 9930
rect 19996 9654 20024 10406
rect 20732 10198 20760 11478
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19536 7002 19564 7142
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 6390 19012 6598
rect 19260 6458 19288 6831
rect 19628 6662 19656 7754
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 6730 19748 7686
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 18972 6384 19024 6390
rect 18972 6326 19024 6332
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19720 5914 19748 6666
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19260 5234 19288 5510
rect 19444 5370 19472 5646
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18432 3534 18460 4490
rect 18524 3942 18552 5034
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18524 3058 18552 3538
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 17972 2746 18184 2774
rect 18248 2746 18368 2774
rect 18156 2378 18184 2746
rect 18340 2530 18368 2746
rect 18248 2502 18368 2530
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18248 800 18276 2502
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18340 1698 18368 2382
rect 18328 1692 18380 1698
rect 18328 1634 18380 1640
rect 18616 800 18644 4966
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19720 4146 19748 4490
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19444 4026 19472 4082
rect 19444 3998 19564 4026
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18984 800 19012 3674
rect 19536 2854 19564 3998
rect 19720 3618 19748 4082
rect 19628 3602 19748 3618
rect 19616 3596 19748 3602
rect 19668 3590 19748 3596
rect 19616 3538 19668 3544
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19352 800 19380 2586
rect 19628 2530 19656 3538
rect 19812 3466 19840 5850
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19536 2502 19656 2530
rect 19536 2446 19564 2502
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19720 800 19748 2586
rect 20088 800 20116 5578
rect 20180 2650 20208 9862
rect 20824 8974 20852 11290
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8090 20668 8774
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20456 5642 20484 6394
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20548 2990 20576 3470
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20732 2774 20760 5510
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20824 3924 20852 5170
rect 20916 4026 20944 9658
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21008 5846 21036 6802
rect 21100 6322 21128 12038
rect 21192 8634 21220 16594
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11762 21404 12038
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21376 11354 21404 11698
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 10674 21404 11290
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21376 10266 21404 10610
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21376 9722 21404 10202
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21376 9042 21404 9658
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21376 8090 21404 8978
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20996 5840 21048 5846
rect 21100 5817 21128 6258
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 20996 5782 21048 5788
rect 21086 5808 21142 5817
rect 21008 5234 21036 5782
rect 21086 5743 21142 5752
rect 21192 5302 21220 6054
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21008 4690 21036 5170
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 21008 4214 21036 4626
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 20916 3998 21036 4026
rect 20824 3896 20944 3924
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20456 2746 20760 2774
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20456 800 20484 2746
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20732 1970 20760 2246
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 20824 800 20852 2994
rect 20916 2310 20944 3896
rect 21008 3534 21036 3998
rect 21100 3738 21128 4422
rect 21284 4146 21312 7958
rect 21376 7546 21404 8026
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21376 7002 21404 7482
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 21468 4622 21496 12174
rect 21560 7313 21588 12650
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21546 7304 21602 7313
rect 21546 7239 21602 7248
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21284 2650 21312 3130
rect 21560 2774 21588 7239
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21468 2746 21588 2774
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21468 2446 21496 2746
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 11716 734 11928 762
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
<< via2 >>
rect 2962 21256 3018 21312
rect 2870 20848 2926 20904
rect 2778 20440 2834 20496
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 1490 18808 1546 18864
rect 1490 18400 1546 18456
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1490 15544 1546 15600
rect 1490 15136 1546 15192
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1490 13912 1546 13968
rect 1490 13504 1546 13560
rect 1490 13096 1546 13152
rect 2042 20052 2098 20088
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 2042 20032 2044 20052
rect 2044 20032 2096 20052
rect 2096 20032 2098 20052
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 2042 19236 2098 19272
rect 2042 19216 2044 19236
rect 2044 19216 2096 19236
rect 2096 19216 2098 19236
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 2042 17584 2098 17640
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 2134 15972 2190 16008
rect 2134 15952 2136 15972
rect 2136 15952 2188 15972
rect 2188 15952 2190 15972
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 2134 14320 2190 14376
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 1398 12688 1454 12744
rect 1490 12280 1546 12336
rect 1214 11736 1270 11792
rect 938 3748 940 3768
rect 940 3748 992 3768
rect 992 3748 994 3768
rect 938 3712 994 3748
rect 1490 11464 1546 11520
rect 1398 10920 1454 10976
rect 1490 10648 1546 10704
rect 1398 10240 1454 10296
rect 1398 9016 1454 9072
rect 1398 8200 1454 8256
rect 1490 8064 1546 8120
rect 1398 7828 1400 7848
rect 1400 7828 1452 7848
rect 1452 7828 1454 7848
rect 1398 7792 1454 7828
rect 1398 6976 1454 7032
rect 1398 6568 1454 6624
rect 1398 6160 1454 6216
rect 1398 5344 1454 5400
rect 1674 10648 1730 10704
rect 1950 11212 2006 11248
rect 1950 11192 1952 11212
rect 1952 11192 2004 11212
rect 2004 11192 2006 11212
rect 1858 9424 1914 9480
rect 1858 8608 1914 8664
rect 2042 9016 2098 9072
rect 2042 8336 2098 8392
rect 1582 6976 1638 7032
rect 1858 7384 1914 7440
rect 1766 6296 1822 6352
rect 1582 5616 1638 5672
rect 1858 4972 1860 4992
rect 1860 4972 1912 4992
rect 1912 4972 1914 4992
rect 1858 4936 1914 4972
rect 1858 4564 1860 4584
rect 1860 4564 1912 4584
rect 1912 4564 1914 4584
rect 1858 4528 1914 4564
rect 2042 7928 2098 7984
rect 2318 9832 2374 9888
rect 2594 11636 2596 11656
rect 2596 11636 2648 11656
rect 2648 11636 2650 11656
rect 2594 11600 2650 11636
rect 2594 10548 2596 10568
rect 2596 10548 2648 10568
rect 2648 10548 2650 10568
rect 2594 10512 2650 10548
rect 2502 9968 2558 10024
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3330 11872 3386 11928
rect 2962 10104 3018 10160
rect 2502 7792 2558 7848
rect 3882 12144 3938 12200
rect 3790 11620 3846 11656
rect 3790 11600 3792 11620
rect 3792 11600 3844 11620
rect 3844 11600 3846 11620
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3054 8064 3110 8120
rect 2870 7520 2926 7576
rect 2226 6860 2282 6896
rect 2226 6840 2228 6860
rect 2228 6840 2280 6860
rect 2280 6840 2282 6860
rect 2318 5072 2374 5128
rect 2226 4140 2282 4176
rect 2226 4120 2228 4140
rect 2228 4120 2280 4140
rect 2280 4120 2282 4140
rect 2042 3576 2098 3632
rect 2962 7268 3018 7304
rect 2962 7248 2964 7268
rect 2964 7248 3016 7268
rect 3016 7248 3018 7268
rect 2778 5752 2834 5808
rect 2778 5208 2834 5264
rect 2778 4936 2834 4992
rect 2778 3032 2834 3088
rect 2962 4936 3018 4992
rect 2962 4528 3018 4584
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3514 9424 3570 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 5722 14320 5778 14376
rect 4066 9832 4122 9888
rect 4066 8608 4122 8664
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4158 8472 4214 8528
rect 3882 6840 3938 6896
rect 2962 2488 3018 2544
rect 4250 7656 4306 7712
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3790 5752 3846 5808
rect 4158 5888 4214 5944
rect 4342 6160 4398 6216
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3606 4664 3662 4720
rect 3974 4120 4030 4176
rect 4526 6024 4582 6080
rect 4986 9696 5042 9752
rect 4986 9424 5042 9480
rect 4802 7384 4858 7440
rect 4434 4256 4490 4312
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3698 3440 3754 3496
rect 3422 3032 3478 3088
rect 3238 2080 3294 2136
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3974 2760 4030 2816
rect 4250 3848 4306 3904
rect 4342 3440 4398 3496
rect 4066 1672 4122 1728
rect 4802 4004 4858 4040
rect 4802 3984 4804 4004
rect 4804 3984 4856 4004
rect 4856 3984 4858 4004
rect 4710 3732 4766 3768
rect 4710 3712 4712 3732
rect 4712 3712 4764 3732
rect 4764 3712 4766 3732
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 5630 11636 5632 11656
rect 5632 11636 5684 11656
rect 5684 11636 5686 11656
rect 5630 11600 5686 11636
rect 5078 4256 5134 4312
rect 6550 11056 6606 11112
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5630 8608 5686 8664
rect 5538 7656 5594 7712
rect 5446 7520 5502 7576
rect 5354 4936 5410 4992
rect 5078 3440 5134 3496
rect 5538 6704 5594 6760
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6734 10784 6790 10840
rect 6734 10512 6790 10568
rect 6918 10532 6974 10568
rect 6918 10512 6920 10532
rect 6920 10512 6972 10532
rect 6972 10512 6974 10532
rect 6550 9560 6606 9616
rect 6642 9424 6698 9480
rect 5906 7112 5962 7168
rect 5906 4664 5962 4720
rect 5722 4256 5778 4312
rect 5446 3984 5502 4040
rect 5630 3848 5686 3904
rect 5538 3188 5594 3224
rect 5538 3168 5540 3188
rect 5540 3168 5592 3188
rect 5592 3168 5594 3188
rect 5906 3848 5962 3904
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 7102 8336 7158 8392
rect 6826 8064 6882 8120
rect 6734 6976 6790 7032
rect 6550 5752 6606 5808
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6734 5092 6790 5128
rect 6734 5072 6736 5092
rect 6736 5072 6788 5092
rect 6788 5072 6790 5092
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6090 3848 6146 3904
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 5998 2916 6054 2952
rect 5998 2896 6000 2916
rect 6000 2896 6052 2916
rect 6052 2896 6054 2916
rect 5906 1808 5962 1864
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 8206 13232 8262 13288
rect 7286 9968 7342 10024
rect 7102 6840 7158 6896
rect 7010 6568 7066 6624
rect 7930 11192 7986 11248
rect 8022 9560 8078 9616
rect 7746 8880 7802 8936
rect 7102 6432 7158 6488
rect 7102 5616 7158 5672
rect 6826 2624 6882 2680
rect 7194 3984 7250 4040
rect 7378 5480 7434 5536
rect 7378 4936 7434 4992
rect 7470 3576 7526 3632
rect 7562 3168 7618 3224
rect 6734 2352 6790 2408
rect 6642 2216 6698 2272
rect 7838 6840 7894 6896
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 9770 13776 9826 13832
rect 10138 13640 10194 13696
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 10230 13232 10286 13288
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9586 12300 9642 12336
rect 9586 12280 9588 12300
rect 9588 12280 9640 12300
rect 9640 12280 9642 12300
rect 9218 11736 9274 11792
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8942 10684 8944 10704
rect 8944 10684 8996 10704
rect 8996 10684 8998 10704
rect 8942 10648 8998 10684
rect 8206 9968 8262 10024
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8206 6976 8262 7032
rect 8022 5752 8078 5808
rect 8206 6160 8262 6216
rect 8114 4392 8170 4448
rect 7838 4120 7894 4176
rect 8298 5788 8300 5808
rect 8300 5788 8352 5808
rect 8352 5788 8354 5808
rect 8298 5752 8354 5788
rect 8298 5344 8354 5400
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8942 7520 8998 7576
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8666 6332 8668 6352
rect 8668 6332 8720 6352
rect 8720 6332 8722 6352
rect 8666 6296 8722 6332
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9402 9696 9458 9752
rect 9770 9016 9826 9072
rect 9954 6604 9956 6624
rect 9956 6604 10008 6624
rect 10008 6604 10010 6624
rect 9954 6568 10010 6604
rect 9678 5480 9734 5536
rect 8482 4936 8538 4992
rect 8114 3440 8170 3496
rect 8114 3032 8170 3088
rect 8390 4120 8446 4176
rect 8298 3576 8354 3632
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9218 4392 9274 4448
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8666 3304 8722 3360
rect 9034 3304 9090 3360
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9310 3576 9366 3632
rect 9494 4528 9550 4584
rect 9494 4256 9550 4312
rect 9770 3984 9826 4040
rect 9494 3712 9550 3768
rect 9310 3304 9366 3360
rect 9494 3188 9550 3224
rect 9494 3168 9496 3188
rect 9496 3168 9548 3188
rect 9548 3168 9550 3188
rect 9218 2624 9274 2680
rect 9770 3168 9826 3224
rect 9678 2488 9734 2544
rect 9954 4972 9956 4992
rect 9956 4972 10008 4992
rect 10008 4972 10010 4992
rect 9954 4936 10010 4972
rect 9954 4004 10010 4040
rect 9954 3984 9956 4004
rect 9956 3984 10008 4004
rect 10008 3984 10010 4004
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11978 13932 12034 13968
rect 11978 13912 11980 13932
rect 11980 13912 12032 13932
rect 12032 13912 12034 13932
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10690 11192 10746 11248
rect 10782 11056 10838 11112
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10138 3032 10194 3088
rect 10874 8336 10930 8392
rect 10690 6432 10746 6488
rect 10782 6160 10838 6216
rect 10966 4528 11022 4584
rect 11794 11328 11850 11384
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11886 8372 11888 8392
rect 11888 8372 11940 8392
rect 11940 8372 11942 8392
rect 11886 8336 11942 8372
rect 11242 7792 11298 7848
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11242 5616 11298 5672
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 10966 2080 11022 2136
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11886 5480 11942 5536
rect 11886 5208 11942 5264
rect 11886 3984 11942 4040
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21270 17176 21326 17232
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 12254 9560 12310 9616
rect 12070 5208 12126 5264
rect 12070 4936 12126 4992
rect 12438 9596 12440 9616
rect 12440 9596 12492 9616
rect 12492 9596 12494 9616
rect 12438 9560 12494 9596
rect 12714 10648 12770 10704
rect 13818 13640 13874 13696
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13450 11600 13506 11656
rect 13266 9968 13322 10024
rect 12070 3848 12126 3904
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12070 1808 12126 1864
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14278 8880 14334 8936
rect 13726 8492 13782 8528
rect 13726 8472 13728 8492
rect 13728 8472 13780 8492
rect 13780 8472 13782 8492
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 15750 9424 15806 9480
rect 15934 10512 15990 10568
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16670 10104 16726 10160
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 17774 10512 17830 10568
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 20534 12180 20536 12200
rect 20536 12180 20588 12200
rect 20588 12180 20590 12200
rect 20534 12144 20590 12180
rect 20810 12280 20866 12336
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 18142 9580 18198 9616
rect 18142 9560 18144 9580
rect 18144 9560 18196 9580
rect 18196 9560 18198 9580
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 17314 8336 17370 8392
rect 15750 6724 15806 6760
rect 15750 6704 15752 6724
rect 15752 6704 15804 6724
rect 15804 6704 15806 6724
rect 15566 5752 15622 5808
rect 14094 5516 14096 5536
rect 14096 5516 14148 5536
rect 14148 5516 14150 5536
rect 14094 5480 14150 5516
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13726 4800 13782 4856
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14278 3612 14280 3632
rect 14280 3612 14332 3632
rect 14332 3612 14334 3632
rect 14278 3576 14334 3612
rect 15842 5616 15898 5672
rect 14554 4528 14610 4584
rect 14370 3440 14426 3496
rect 13358 2932 13360 2952
rect 13360 2932 13412 2952
rect 13412 2932 13414 2952
rect 13358 2896 13414 2932
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16946 5208 17002 5264
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 15198 1944 15254 2000
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17130 3984 17186 4040
rect 15934 2352 15990 2408
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 18510 7964 18512 7984
rect 18512 7964 18564 7984
rect 18564 7964 18566 7984
rect 18510 7928 18566 7964
rect 17958 7384 18014 7440
rect 18142 5072 18198 5128
rect 18050 4120 18106 4176
rect 17222 3032 17278 3088
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19246 6840 19302 6896
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21086 5752 21142 5808
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21546 7248 21602 7304
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21314 800 21344
rect 2957 21314 3023 21317
rect 0 21312 3023 21314
rect 0 21256 2962 21312
rect 3018 21256 3023 21312
rect 0 21254 3023 21256
rect 0 21224 800 21254
rect 2957 21251 3023 21254
rect 0 20906 800 20936
rect 2865 20906 2931 20909
rect 0 20904 2931 20906
rect 0 20848 2870 20904
rect 2926 20848 2931 20904
rect 0 20846 2931 20848
rect 0 20816 800 20846
rect 2865 20843 2931 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 2773 20498 2839 20501
rect 0 20496 2839 20498
rect 0 20440 2778 20496
rect 2834 20440 2839 20496
rect 0 20438 2839 20440
rect 0 20408 800 20438
rect 2773 20435 2839 20438
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 2037 20090 2103 20093
rect 0 20088 2103 20090
rect 0 20032 2042 20088
rect 2098 20032 2103 20088
rect 0 20030 2103 20032
rect 0 20000 800 20030
rect 2037 20027 2103 20030
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 0 19274 800 19304
rect 2037 19274 2103 19277
rect 0 19272 2103 19274
rect 0 19216 2042 19272
rect 2098 19216 2103 19272
rect 0 19214 2103 19216
rect 0 19184 800 19214
rect 2037 19211 2103 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 0 17642 800 17672
rect 2037 17642 2103 17645
rect 0 17640 2103 17642
rect 0 17584 2042 17640
rect 2098 17584 2103 17640
rect 0 17582 2103 17584
rect 0 17552 800 17582
rect 2037 17579 2103 17582
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 21265 17234 21331 17237
rect 22200 17234 23000 17264
rect 21265 17232 23000 17234
rect 21265 17176 21270 17232
rect 21326 17176 23000 17232
rect 21265 17174 23000 17176
rect 21265 17171 21331 17174
rect 22200 17144 23000 17174
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 0 16010 800 16040
rect 2129 16010 2195 16013
rect 0 16008 2195 16010
rect 0 15952 2134 16008
rect 2190 15952 2195 16008
rect 0 15950 2195 15952
rect 0 15920 800 15950
rect 2129 15947 2195 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 0 14378 800 14408
rect 2129 14378 2195 14381
rect 0 14376 2195 14378
rect 0 14320 2134 14376
rect 2190 14320 2195 14376
rect 0 14318 2195 14320
rect 0 14288 800 14318
rect 2129 14315 2195 14318
rect 5717 14378 5783 14381
rect 9990 14378 9996 14380
rect 5717 14376 9996 14378
rect 5717 14320 5722 14376
rect 5778 14320 9996 14376
rect 5717 14318 9996 14320
rect 5717 14315 5783 14318
rect 9990 14316 9996 14318
rect 10060 14316 10066 14380
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 0 13970 800 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 800 13910
rect 1485 13907 1551 13910
rect 9438 13908 9444 13972
rect 9508 13970 9514 13972
rect 11973 13970 12039 13973
rect 9508 13968 12039 13970
rect 9508 13912 11978 13968
rect 12034 13912 12039 13968
rect 9508 13910 12039 13912
rect 9508 13908 9514 13910
rect 11973 13907 12039 13910
rect 9765 13836 9831 13837
rect 9765 13832 9812 13836
rect 9876 13834 9882 13836
rect 9765 13776 9770 13832
rect 9765 13772 9812 13776
rect 9876 13774 9922 13834
rect 9876 13772 9882 13774
rect 9765 13771 9831 13772
rect 10133 13698 10199 13701
rect 13813 13698 13879 13701
rect 10133 13696 13879 13698
rect 10133 13640 10138 13696
rect 10194 13640 13818 13696
rect 13874 13640 13879 13696
rect 10133 13638 13879 13640
rect 10133 13635 10199 13638
rect 13813 13635 13879 13638
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 1485 13562 1551 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 8201 13290 8267 13293
rect 10225 13290 10291 13293
rect 8201 13288 10291 13290
rect 8201 13232 8206 13288
rect 8262 13232 10230 13288
rect 10286 13232 10291 13288
rect 8201 13230 10291 13232
rect 8201 13227 8267 13230
rect 10225 13227 10291 13230
rect 0 13154 800 13184
rect 1485 13154 1551 13157
rect 0 13152 1551 13154
rect 0 13096 1490 13152
rect 1546 13096 1551 13152
rect 0 13094 1551 13096
rect 0 13064 800 13094
rect 1485 13091 1551 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 0 12746 800 12776
rect 1393 12746 1459 12749
rect 0 12744 1459 12746
rect 0 12688 1398 12744
rect 1454 12688 1459 12744
rect 0 12686 1459 12688
rect 0 12656 800 12686
rect 1393 12683 1459 12686
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 9581 12338 9647 12341
rect 20805 12338 20871 12341
rect 9581 12336 20871 12338
rect 9581 12280 9586 12336
rect 9642 12280 20810 12336
rect 20866 12280 20871 12336
rect 9581 12278 20871 12280
rect 9581 12275 9647 12278
rect 20805 12275 20871 12278
rect 3877 12202 3943 12205
rect 20529 12202 20595 12205
rect 3877 12200 20595 12202
rect 3877 12144 3882 12200
rect 3938 12144 20534 12200
rect 20590 12144 20595 12200
rect 3877 12142 20595 12144
rect 3877 12139 3943 12142
rect 20529 12139 20595 12142
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 3325 11930 3391 11933
rect 0 11928 3391 11930
rect 0 11872 3330 11928
rect 3386 11872 3391 11928
rect 0 11870 3391 11872
rect 0 11840 800 11870
rect 3325 11867 3391 11870
rect 1209 11794 1275 11797
rect 9213 11794 9279 11797
rect 1209 11792 9279 11794
rect 1209 11736 1214 11792
rect 1270 11736 9218 11792
rect 9274 11736 9279 11792
rect 1209 11734 9279 11736
rect 1209 11731 1275 11734
rect 9213 11731 9279 11734
rect 2589 11658 2655 11661
rect 3785 11658 3851 11661
rect 2589 11656 3851 11658
rect 2589 11600 2594 11656
rect 2650 11600 3790 11656
rect 3846 11600 3851 11656
rect 2589 11598 3851 11600
rect 2589 11595 2655 11598
rect 3785 11595 3851 11598
rect 5625 11658 5691 11661
rect 13445 11658 13511 11661
rect 5625 11656 13511 11658
rect 5625 11600 5630 11656
rect 5686 11600 13450 11656
rect 13506 11600 13511 11656
rect 5625 11598 13511 11600
rect 5625 11595 5691 11598
rect 13445 11595 13511 11598
rect 0 11522 800 11552
rect 1485 11522 1551 11525
rect 0 11520 1551 11522
rect 0 11464 1490 11520
rect 1546 11464 1551 11520
rect 0 11462 1551 11464
rect 0 11432 800 11462
rect 1485 11459 1551 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 11789 11386 11855 11389
rect 5398 11326 8586 11386
rect 1945 11250 2011 11253
rect 5398 11250 5458 11326
rect 1945 11248 5458 11250
rect 1945 11192 1950 11248
rect 2006 11192 5458 11248
rect 1945 11190 5458 11192
rect 1945 11187 2011 11190
rect 5574 11188 5580 11252
rect 5644 11250 5650 11252
rect 7925 11250 7991 11253
rect 5644 11248 7991 11250
rect 5644 11192 7930 11248
rect 7986 11192 7991 11248
rect 5644 11190 7991 11192
rect 8526 11250 8586 11326
rect 9446 11384 11855 11386
rect 9446 11328 11794 11384
rect 11850 11328 11855 11384
rect 9446 11326 11855 11328
rect 9446 11250 9506 11326
rect 11789 11323 11855 11326
rect 8526 11190 9506 11250
rect 5644 11188 5650 11190
rect 7925 11187 7991 11190
rect 9622 11188 9628 11252
rect 9692 11250 9698 11252
rect 10685 11250 10751 11253
rect 9692 11248 10751 11250
rect 9692 11192 10690 11248
rect 10746 11192 10751 11248
rect 9692 11190 10751 11192
rect 9692 11188 9698 11190
rect 10685 11187 10751 11190
rect 0 11114 800 11144
rect 6545 11114 6611 11117
rect 6678 11114 6684 11116
rect 0 11054 1456 11114
rect 0 11024 800 11054
rect 1396 10981 1456 11054
rect 6545 11112 6684 11114
rect 6545 11056 6550 11112
rect 6606 11056 6684 11112
rect 6545 11054 6684 11056
rect 6545 11051 6611 11054
rect 6678 11052 6684 11054
rect 6748 11052 6754 11116
rect 10777 11114 10843 11117
rect 10910 11114 10916 11116
rect 10777 11112 10916 11114
rect 10777 11056 10782 11112
rect 10838 11056 10916 11112
rect 10777 11054 10916 11056
rect 10777 11051 10843 11054
rect 10910 11052 10916 11054
rect 10980 11052 10986 11116
rect 1393 10976 1459 10981
rect 1393 10920 1398 10976
rect 1454 10920 1459 10976
rect 1393 10915 1459 10920
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 6729 10842 6795 10845
rect 6729 10840 9690 10842
rect 6729 10784 6734 10840
rect 6790 10784 9690 10840
rect 6729 10782 9690 10784
rect 6729 10779 6795 10782
rect 0 10706 800 10736
rect 1485 10706 1551 10709
rect 0 10704 1551 10706
rect 0 10648 1490 10704
rect 1546 10648 1551 10704
rect 0 10646 1551 10648
rect 0 10616 800 10646
rect 1485 10643 1551 10646
rect 1669 10706 1735 10709
rect 8937 10706 9003 10709
rect 1669 10704 9003 10706
rect 1669 10648 1674 10704
rect 1730 10648 8942 10704
rect 8998 10648 9003 10704
rect 1669 10646 9003 10648
rect 9630 10706 9690 10782
rect 12709 10706 12775 10709
rect 9630 10704 12775 10706
rect 9630 10648 12714 10704
rect 12770 10648 12775 10704
rect 9630 10646 12775 10648
rect 1669 10643 1735 10646
rect 8937 10643 9003 10646
rect 12709 10643 12775 10646
rect 2589 10570 2655 10573
rect 6729 10570 6795 10573
rect 2589 10568 6795 10570
rect 2589 10512 2594 10568
rect 2650 10512 6734 10568
rect 6790 10512 6795 10568
rect 2589 10510 6795 10512
rect 2589 10507 2655 10510
rect 6729 10507 6795 10510
rect 6913 10570 6979 10573
rect 15929 10570 15995 10573
rect 17769 10570 17835 10573
rect 6913 10568 17835 10570
rect 6913 10512 6918 10568
rect 6974 10512 15934 10568
rect 15990 10512 17774 10568
rect 17830 10512 17835 10568
rect 6913 10510 17835 10512
rect 6913 10507 6979 10510
rect 15929 10507 15995 10510
rect 17769 10507 17835 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 2957 10162 3023 10165
rect 16665 10162 16731 10165
rect 2957 10160 16731 10162
rect 2957 10104 2962 10160
rect 3018 10104 16670 10160
rect 16726 10104 16731 10160
rect 2957 10102 16731 10104
rect 2957 10099 3023 10102
rect 16665 10099 16731 10102
rect 2497 10026 2563 10029
rect 7281 10026 7347 10029
rect 2497 10024 7347 10026
rect 2497 9968 2502 10024
rect 2558 9968 7286 10024
rect 7342 9968 7347 10024
rect 2497 9966 7347 9968
rect 2497 9963 2563 9966
rect 7281 9963 7347 9966
rect 8201 10026 8267 10029
rect 13261 10026 13327 10029
rect 8201 10024 13327 10026
rect 8201 9968 8206 10024
rect 8262 9968 13266 10024
rect 13322 9968 13327 10024
rect 8201 9966 13327 9968
rect 8201 9963 8267 9966
rect 13261 9963 13327 9966
rect 0 9890 800 9920
rect 2313 9890 2379 9893
rect 0 9888 2379 9890
rect 0 9832 2318 9888
rect 2374 9832 2379 9888
rect 0 9830 2379 9832
rect 0 9800 800 9830
rect 2313 9827 2379 9830
rect 3918 9828 3924 9892
rect 3988 9890 3994 9892
rect 4061 9890 4127 9893
rect 3988 9888 4127 9890
rect 3988 9832 4066 9888
rect 4122 9832 4127 9888
rect 3988 9830 4127 9832
rect 3988 9828 3994 9830
rect 4061 9827 4127 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 4470 9692 4476 9756
rect 4540 9754 4546 9756
rect 4981 9754 5047 9757
rect 4540 9752 5047 9754
rect 4540 9696 4986 9752
rect 5042 9696 5047 9752
rect 4540 9694 5047 9696
rect 4540 9692 4546 9694
rect 4981 9691 5047 9694
rect 8150 9692 8156 9756
rect 8220 9754 8226 9756
rect 9397 9754 9463 9757
rect 8220 9752 9463 9754
rect 8220 9696 9402 9752
rect 9458 9696 9463 9752
rect 8220 9694 9463 9696
rect 8220 9692 8226 9694
rect 9397 9691 9463 9694
rect 2814 9556 2820 9620
rect 2884 9618 2890 9620
rect 6545 9618 6611 9621
rect 2884 9616 6611 9618
rect 2884 9560 6550 9616
rect 6606 9560 6611 9616
rect 2884 9558 6611 9560
rect 2884 9556 2890 9558
rect 6545 9555 6611 9558
rect 8017 9618 8083 9621
rect 12249 9618 12315 9621
rect 8017 9616 12315 9618
rect 8017 9560 8022 9616
rect 8078 9560 12254 9616
rect 12310 9560 12315 9616
rect 8017 9558 12315 9560
rect 8017 9555 8083 9558
rect 12249 9555 12315 9558
rect 12433 9618 12499 9621
rect 18137 9618 18203 9621
rect 12433 9616 18203 9618
rect 12433 9560 12438 9616
rect 12494 9560 18142 9616
rect 18198 9560 18203 9616
rect 12433 9558 18203 9560
rect 12433 9555 12499 9558
rect 18137 9555 18203 9558
rect 0 9482 800 9512
rect 1853 9482 1919 9485
rect 0 9480 1919 9482
rect 0 9424 1858 9480
rect 1914 9424 1919 9480
rect 0 9422 1919 9424
rect 0 9392 800 9422
rect 1853 9419 1919 9422
rect 3366 9420 3372 9484
rect 3436 9482 3442 9484
rect 3509 9482 3575 9485
rect 3436 9480 3575 9482
rect 3436 9424 3514 9480
rect 3570 9424 3575 9480
rect 3436 9422 3575 9424
rect 3436 9420 3442 9422
rect 3509 9419 3575 9422
rect 4654 9420 4660 9484
rect 4724 9482 4730 9484
rect 4981 9482 5047 9485
rect 4724 9480 5047 9482
rect 4724 9424 4986 9480
rect 5042 9424 5047 9480
rect 4724 9422 5047 9424
rect 4724 9420 4730 9422
rect 4981 9419 5047 9422
rect 6637 9482 6703 9485
rect 15745 9482 15811 9485
rect 6637 9480 15811 9482
rect 6637 9424 6642 9480
rect 6698 9424 15750 9480
rect 15806 9424 15811 9480
rect 6637 9422 15811 9424
rect 6637 9419 6703 9422
rect 15745 9419 15811 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 2037 9074 2103 9077
rect 9765 9074 9831 9077
rect 2037 9072 9831 9074
rect 2037 9016 2042 9072
rect 2098 9016 9770 9072
rect 9826 9016 9831 9072
rect 2037 9014 9831 9016
rect 2037 9011 2103 9014
rect 9765 9011 9831 9014
rect 7741 8938 7807 8941
rect 14273 8938 14339 8941
rect 7741 8936 14339 8938
rect 7741 8880 7746 8936
rect 7802 8880 14278 8936
rect 14334 8880 14339 8936
rect 7741 8878 14339 8880
rect 7741 8875 7807 8878
rect 14273 8875 14339 8878
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 1853 8666 1919 8669
rect 0 8664 1919 8666
rect 0 8608 1858 8664
rect 1914 8608 1919 8664
rect 0 8606 1919 8608
rect 0 8576 800 8606
rect 1853 8603 1919 8606
rect 4061 8668 4127 8669
rect 4061 8664 4108 8668
rect 4172 8666 4178 8668
rect 4061 8608 4066 8664
rect 4061 8604 4108 8608
rect 4172 8606 4218 8666
rect 4172 8604 4178 8606
rect 4286 8604 4292 8668
rect 4356 8666 4362 8668
rect 5625 8666 5691 8669
rect 4356 8664 5691 8666
rect 4356 8608 5630 8664
rect 5686 8608 5691 8664
rect 4356 8606 5691 8608
rect 4356 8604 4362 8606
rect 4061 8603 4127 8604
rect 5625 8603 5691 8606
rect 4153 8530 4219 8533
rect 13721 8530 13787 8533
rect 4153 8528 13787 8530
rect 4153 8472 4158 8528
rect 4214 8472 13726 8528
rect 13782 8472 13787 8528
rect 4153 8470 13787 8472
rect 4153 8467 4219 8470
rect 13721 8467 13787 8470
rect 2037 8394 2103 8397
rect 2262 8394 2268 8396
rect 2037 8392 2268 8394
rect 2037 8336 2042 8392
rect 2098 8336 2268 8392
rect 2037 8334 2268 8336
rect 2037 8331 2103 8334
rect 2262 8332 2268 8334
rect 2332 8332 2338 8396
rect 5022 8332 5028 8396
rect 5092 8394 5098 8396
rect 7097 8394 7163 8397
rect 5092 8392 7163 8394
rect 5092 8336 7102 8392
rect 7158 8336 7163 8392
rect 5092 8334 7163 8336
rect 5092 8332 5098 8334
rect 7097 8331 7163 8334
rect 10174 8332 10180 8396
rect 10244 8394 10250 8396
rect 10869 8394 10935 8397
rect 10244 8392 10935 8394
rect 10244 8336 10874 8392
rect 10930 8336 10935 8392
rect 10244 8334 10935 8336
rect 10244 8332 10250 8334
rect 10869 8331 10935 8334
rect 11881 8394 11947 8397
rect 17309 8394 17375 8397
rect 11881 8392 17375 8394
rect 11881 8336 11886 8392
rect 11942 8336 17314 8392
rect 17370 8336 17375 8392
rect 11881 8334 17375 8336
rect 11881 8331 11947 8334
rect 17309 8331 17375 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 1485 8122 1551 8125
rect 3049 8122 3115 8125
rect 1485 8120 3115 8122
rect 1485 8064 1490 8120
rect 1546 8064 3054 8120
rect 3110 8064 3115 8120
rect 1485 8062 3115 8064
rect 1485 8059 1551 8062
rect 3049 8059 3115 8062
rect 6821 8124 6887 8125
rect 6821 8120 6868 8124
rect 6932 8122 6938 8124
rect 6821 8064 6826 8120
rect 6821 8060 6868 8064
rect 6932 8062 6978 8122
rect 6932 8060 6938 8062
rect 6821 8059 6887 8060
rect 2037 7986 2103 7989
rect 18505 7986 18571 7989
rect 2037 7984 18571 7986
rect 2037 7928 2042 7984
rect 2098 7928 18510 7984
rect 18566 7928 18571 7984
rect 2037 7926 18571 7928
rect 2037 7923 2103 7926
rect 18505 7923 18571 7926
rect 0 7850 800 7880
rect 1393 7850 1459 7853
rect 0 7848 1459 7850
rect 0 7792 1398 7848
rect 1454 7792 1459 7848
rect 0 7790 1459 7792
rect 0 7760 800 7790
rect 1393 7787 1459 7790
rect 2497 7850 2563 7853
rect 11237 7850 11303 7853
rect 2497 7848 11303 7850
rect 2497 7792 2502 7848
rect 2558 7792 11242 7848
rect 11298 7792 11303 7848
rect 2497 7790 11303 7792
rect 2497 7787 2563 7790
rect 11237 7787 11303 7790
rect 4245 7714 4311 7717
rect 5533 7714 5599 7717
rect 4245 7712 5599 7714
rect 4245 7656 4250 7712
rect 4306 7656 5538 7712
rect 5594 7656 5599 7712
rect 4245 7654 5599 7656
rect 4245 7651 4311 7654
rect 5533 7651 5599 7654
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 2865 7578 2931 7581
rect 5441 7578 5507 7581
rect 2865 7576 5507 7578
rect 2865 7520 2870 7576
rect 2926 7520 5446 7576
rect 5502 7520 5507 7576
rect 2865 7518 5507 7520
rect 2865 7515 2931 7518
rect 5441 7515 5507 7518
rect 8334 7516 8340 7580
rect 8404 7578 8410 7580
rect 8937 7578 9003 7581
rect 8404 7576 9003 7578
rect 8404 7520 8942 7576
rect 8998 7520 9003 7576
rect 8404 7518 9003 7520
rect 8404 7516 8410 7518
rect 8937 7515 9003 7518
rect 0 7442 800 7472
rect 1853 7442 1919 7445
rect 0 7440 1919 7442
rect 0 7384 1858 7440
rect 1914 7384 1919 7440
rect 0 7382 1919 7384
rect 0 7352 800 7382
rect 1853 7379 1919 7382
rect 4797 7442 4863 7445
rect 17953 7442 18019 7445
rect 4797 7440 18019 7442
rect 4797 7384 4802 7440
rect 4858 7384 17958 7440
rect 18014 7384 18019 7440
rect 4797 7382 18019 7384
rect 4797 7379 4863 7382
rect 17953 7379 18019 7382
rect 2957 7306 3023 7309
rect 21541 7306 21607 7309
rect 2957 7304 21607 7306
rect 2957 7248 2962 7304
rect 3018 7248 21546 7304
rect 21602 7248 21607 7304
rect 2957 7246 21607 7248
rect 2957 7243 3023 7246
rect 21541 7243 21607 7246
rect 5758 7108 5764 7172
rect 5828 7170 5834 7172
rect 5901 7170 5967 7173
rect 5828 7168 5967 7170
rect 5828 7112 5906 7168
rect 5962 7112 5967 7168
rect 5828 7110 5967 7112
rect 5828 7108 5834 7110
rect 5901 7107 5967 7110
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 1393 7034 1459 7037
rect 0 7032 1459 7034
rect 0 6976 1398 7032
rect 1454 6976 1459 7032
rect 0 6974 1459 6976
rect 0 6944 800 6974
rect 1393 6971 1459 6974
rect 1577 7034 1643 7037
rect 2446 7034 2452 7036
rect 1577 7032 2452 7034
rect 1577 6976 1582 7032
rect 1638 6976 2452 7032
rect 1577 6974 2452 6976
rect 1577 6971 1643 6974
rect 2446 6972 2452 6974
rect 2516 6972 2522 7036
rect 4838 6972 4844 7036
rect 4908 7034 4914 7036
rect 6729 7034 6795 7037
rect 4908 7032 6795 7034
rect 4908 6976 6734 7032
rect 6790 6976 6795 7032
rect 4908 6974 6795 6976
rect 4908 6972 4914 6974
rect 6729 6971 6795 6974
rect 7230 6972 7236 7036
rect 7300 7034 7306 7036
rect 8201 7034 8267 7037
rect 7300 7032 8267 7034
rect 7300 6976 8206 7032
rect 8262 6976 8267 7032
rect 7300 6974 8267 6976
rect 7300 6972 7306 6974
rect 8201 6971 8267 6974
rect 2221 6898 2287 6901
rect 3877 6898 3943 6901
rect 7097 6898 7163 6901
rect 2221 6896 7163 6898
rect 2221 6840 2226 6896
rect 2282 6840 3882 6896
rect 3938 6840 7102 6896
rect 7158 6840 7163 6896
rect 2221 6838 7163 6840
rect 2221 6835 2287 6838
rect 3877 6835 3943 6838
rect 7097 6835 7163 6838
rect 7833 6898 7899 6901
rect 19241 6898 19307 6901
rect 7833 6896 19307 6898
rect 7833 6840 7838 6896
rect 7894 6840 19246 6896
rect 19302 6840 19307 6896
rect 7833 6838 19307 6840
rect 7833 6835 7899 6838
rect 19241 6835 19307 6838
rect 5533 6762 5599 6765
rect 15745 6762 15811 6765
rect 5533 6760 15811 6762
rect 5533 6704 5538 6760
rect 5594 6704 15750 6760
rect 15806 6704 15811 6760
rect 5533 6702 15811 6704
rect 5533 6699 5599 6702
rect 15745 6699 15811 6702
rect 0 6626 800 6656
rect 1393 6626 1459 6629
rect 0 6624 1459 6626
rect 0 6568 1398 6624
rect 1454 6568 1459 6624
rect 0 6566 1459 6568
rect 0 6536 800 6566
rect 1393 6563 1459 6566
rect 7005 6626 7071 6629
rect 9949 6626 10015 6629
rect 7005 6624 10015 6626
rect 7005 6568 7010 6624
rect 7066 6568 9954 6624
rect 10010 6568 10015 6624
rect 7005 6566 10015 6568
rect 7005 6563 7071 6566
rect 9949 6563 10015 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 7097 6490 7163 6493
rect 10685 6490 10751 6493
rect 7097 6488 10751 6490
rect 7097 6432 7102 6488
rect 7158 6432 10690 6488
rect 10746 6432 10751 6488
rect 7097 6430 10751 6432
rect 7097 6427 7163 6430
rect 10685 6427 10751 6430
rect 1761 6354 1827 6357
rect 8661 6354 8727 6357
rect 1761 6352 8727 6354
rect 1761 6296 1766 6352
rect 1822 6296 8666 6352
rect 8722 6296 8727 6352
rect 1761 6294 8727 6296
rect 1761 6291 1827 6294
rect 8661 6291 8727 6294
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 4337 6218 4403 6221
rect 8201 6218 8267 6221
rect 10777 6218 10843 6221
rect 4337 6216 8267 6218
rect 4337 6160 4342 6216
rect 4398 6160 8206 6216
rect 8262 6160 8267 6216
rect 4337 6158 8267 6160
rect 4337 6155 4403 6158
rect 8201 6155 8267 6158
rect 8526 6216 10843 6218
rect 8526 6160 10782 6216
rect 10838 6160 10843 6216
rect 8526 6158 10843 6160
rect 4521 6082 4587 6085
rect 8526 6082 8586 6158
rect 10777 6155 10843 6158
rect 4521 6080 8586 6082
rect 4521 6024 4526 6080
rect 4582 6024 8586 6080
rect 4521 6022 8586 6024
rect 4521 6019 4587 6022
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 4153 5946 4219 5949
rect 7414 5946 7420 5948
rect 4153 5944 7420 5946
rect 4153 5888 4158 5944
rect 4214 5888 7420 5944
rect 4153 5886 7420 5888
rect 4153 5883 4219 5886
rect 7414 5884 7420 5886
rect 7484 5884 7490 5948
rect 0 5810 800 5840
rect 2773 5810 2839 5813
rect 0 5808 2839 5810
rect 0 5752 2778 5808
rect 2834 5752 2839 5808
rect 0 5750 2839 5752
rect 0 5720 800 5750
rect 2773 5747 2839 5750
rect 3785 5810 3851 5813
rect 6545 5810 6611 5813
rect 3785 5808 6611 5810
rect 3785 5752 3790 5808
rect 3846 5752 6550 5808
rect 6606 5752 6611 5808
rect 3785 5750 6611 5752
rect 3785 5747 3851 5750
rect 6545 5747 6611 5750
rect 7046 5748 7052 5812
rect 7116 5810 7122 5812
rect 8017 5810 8083 5813
rect 7116 5808 8083 5810
rect 7116 5752 8022 5808
rect 8078 5752 8083 5808
rect 7116 5750 8083 5752
rect 7116 5748 7122 5750
rect 8017 5747 8083 5750
rect 8293 5810 8359 5813
rect 15561 5810 15627 5813
rect 8293 5808 15627 5810
rect 8293 5752 8298 5808
rect 8354 5752 15566 5808
rect 15622 5752 15627 5808
rect 8293 5750 15627 5752
rect 8293 5747 8359 5750
rect 15561 5747 15627 5750
rect 21081 5810 21147 5813
rect 22200 5810 23000 5840
rect 21081 5808 23000 5810
rect 21081 5752 21086 5808
rect 21142 5752 23000 5808
rect 21081 5750 23000 5752
rect 21081 5747 21147 5750
rect 22200 5720 23000 5750
rect 1577 5674 1643 5677
rect 7097 5674 7163 5677
rect 1577 5672 7163 5674
rect 1577 5616 1582 5672
rect 1638 5616 7102 5672
rect 7158 5616 7163 5672
rect 1577 5614 7163 5616
rect 1577 5611 1643 5614
rect 7097 5611 7163 5614
rect 11237 5674 11303 5677
rect 15837 5674 15903 5677
rect 11237 5672 15903 5674
rect 11237 5616 11242 5672
rect 11298 5616 15842 5672
rect 15898 5616 15903 5672
rect 11237 5614 15903 5616
rect 11237 5611 11303 5614
rect 15837 5611 15903 5614
rect 7373 5538 7439 5541
rect 9673 5538 9739 5541
rect 7373 5536 9739 5538
rect 7373 5480 7378 5536
rect 7434 5480 9678 5536
rect 9734 5480 9739 5536
rect 7373 5478 9739 5480
rect 7373 5475 7439 5478
rect 9673 5475 9739 5478
rect 11881 5538 11947 5541
rect 14089 5538 14155 5541
rect 11881 5536 14155 5538
rect 11881 5480 11886 5536
rect 11942 5480 14094 5536
rect 14150 5480 14155 5536
rect 11881 5478 14155 5480
rect 11881 5475 11947 5478
rect 14089 5475 14155 5478
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 1393 5402 1459 5405
rect 0 5400 1459 5402
rect 0 5344 1398 5400
rect 1454 5344 1459 5400
rect 0 5342 1459 5344
rect 0 5312 800 5342
rect 1393 5339 1459 5342
rect 7598 5340 7604 5404
rect 7668 5402 7674 5404
rect 8293 5402 8359 5405
rect 7668 5400 8359 5402
rect 7668 5344 8298 5400
rect 8354 5344 8359 5400
rect 7668 5342 8359 5344
rect 7668 5340 7674 5342
rect 8293 5339 8359 5342
rect 2773 5266 2839 5269
rect 11881 5266 11947 5269
rect 2773 5264 11947 5266
rect 2773 5208 2778 5264
rect 2834 5208 11886 5264
rect 11942 5208 11947 5264
rect 2773 5206 11947 5208
rect 2773 5203 2839 5206
rect 11881 5203 11947 5206
rect 12065 5266 12131 5269
rect 16941 5266 17007 5269
rect 12065 5264 17007 5266
rect 12065 5208 12070 5264
rect 12126 5208 16946 5264
rect 17002 5208 17007 5264
rect 12065 5206 17007 5208
rect 12065 5203 12131 5206
rect 16941 5203 17007 5206
rect 2313 5130 2379 5133
rect 6729 5130 6795 5133
rect 18137 5130 18203 5133
rect 2313 5128 5274 5130
rect 2313 5072 2318 5128
rect 2374 5072 5274 5128
rect 2313 5070 5274 5072
rect 2313 5067 2379 5070
rect 0 4994 800 5024
rect 1853 4994 1919 4997
rect 0 4992 1919 4994
rect 0 4936 1858 4992
rect 1914 4936 1919 4992
rect 0 4934 1919 4936
rect 0 4904 800 4934
rect 1853 4931 1919 4934
rect 2773 4994 2839 4997
rect 2957 4994 3023 4997
rect 2773 4992 3023 4994
rect 2773 4936 2778 4992
rect 2834 4936 2962 4992
rect 3018 4936 3023 4992
rect 2773 4934 3023 4936
rect 2773 4931 2839 4934
rect 2957 4931 3023 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 5214 4858 5274 5070
rect 6729 5128 18203 5130
rect 6729 5072 6734 5128
rect 6790 5072 18142 5128
rect 18198 5072 18203 5128
rect 6729 5070 18203 5072
rect 6729 5067 6795 5070
rect 18137 5067 18203 5070
rect 5349 4994 5415 4997
rect 5942 4994 5948 4996
rect 5349 4992 5948 4994
rect 5349 4936 5354 4992
rect 5410 4936 5948 4992
rect 5349 4934 5948 4936
rect 5349 4931 5415 4934
rect 5942 4932 5948 4934
rect 6012 4994 6018 4996
rect 7373 4994 7439 4997
rect 8477 4994 8543 4997
rect 6012 4992 7439 4994
rect 6012 4936 7378 4992
rect 7434 4936 7439 4992
rect 6012 4934 7439 4936
rect 6012 4932 6018 4934
rect 7373 4931 7439 4934
rect 7606 4992 8543 4994
rect 7606 4936 8482 4992
rect 8538 4936 8543 4992
rect 7606 4934 8543 4936
rect 7606 4858 7666 4934
rect 8477 4931 8543 4934
rect 9949 4994 10015 4997
rect 12065 4994 12131 4997
rect 9949 4992 12131 4994
rect 9949 4936 9954 4992
rect 10010 4936 12070 4992
rect 12126 4936 12131 4992
rect 9949 4934 12131 4936
rect 9949 4931 10015 4934
rect 12065 4931 12131 4934
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 13721 4858 13787 4861
rect 5214 4798 7666 4858
rect 12390 4856 13787 4858
rect 12390 4800 13726 4856
rect 13782 4800 13787 4856
rect 12390 4798 13787 4800
rect 3601 4722 3667 4725
rect 3918 4722 3924 4724
rect 3601 4720 3924 4722
rect 3601 4664 3606 4720
rect 3662 4664 3924 4720
rect 3601 4662 3924 4664
rect 3601 4659 3667 4662
rect 3918 4660 3924 4662
rect 3988 4660 3994 4724
rect 5901 4722 5967 4725
rect 12390 4722 12450 4798
rect 13721 4795 13787 4798
rect 5901 4720 12450 4722
rect 5901 4664 5906 4720
rect 5962 4664 12450 4720
rect 5901 4662 12450 4664
rect 5901 4659 5967 4662
rect 0 4586 800 4616
rect 1853 4586 1919 4589
rect 0 4584 1919 4586
rect 0 4528 1858 4584
rect 1914 4528 1919 4584
rect 0 4526 1919 4528
rect 0 4496 800 4526
rect 1853 4523 1919 4526
rect 2957 4586 3023 4589
rect 5758 4586 5764 4588
rect 2957 4584 5764 4586
rect 2957 4528 2962 4584
rect 3018 4528 5764 4584
rect 2957 4526 5764 4528
rect 2957 4523 3023 4526
rect 5758 4524 5764 4526
rect 5828 4524 5834 4588
rect 9489 4586 9555 4589
rect 5950 4584 9555 4586
rect 5950 4528 9494 4584
rect 9550 4528 9555 4584
rect 5950 4526 9555 4528
rect 2262 4388 2268 4452
rect 2332 4450 2338 4452
rect 5950 4450 6010 4526
rect 9489 4523 9555 4526
rect 10961 4586 11027 4589
rect 14549 4586 14615 4589
rect 10961 4584 14615 4586
rect 10961 4528 10966 4584
rect 11022 4528 14554 4584
rect 14610 4528 14615 4584
rect 10961 4526 14615 4528
rect 10961 4523 11027 4526
rect 14549 4523 14615 4526
rect 2332 4390 6010 4450
rect 8109 4450 8175 4453
rect 9213 4450 9279 4453
rect 8109 4448 9279 4450
rect 8109 4392 8114 4448
rect 8170 4392 9218 4448
rect 9274 4392 9279 4448
rect 8109 4390 9279 4392
rect 2332 4388 2338 4390
rect 8109 4387 8175 4390
rect 9213 4387 9279 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 4429 4316 4495 4317
rect 4429 4314 4476 4316
rect 4384 4312 4476 4314
rect 4384 4256 4434 4312
rect 4384 4254 4476 4256
rect 4429 4252 4476 4254
rect 4540 4252 4546 4316
rect 5073 4314 5139 4317
rect 5717 4314 5783 4317
rect 5073 4312 5783 4314
rect 5073 4256 5078 4312
rect 5134 4256 5722 4312
rect 5778 4256 5783 4312
rect 5073 4254 5783 4256
rect 4429 4251 4495 4252
rect 5073 4251 5139 4254
rect 5717 4251 5783 4254
rect 7782 4252 7788 4316
rect 7852 4314 7858 4316
rect 9489 4314 9555 4317
rect 7852 4312 9555 4314
rect 7852 4256 9494 4312
rect 9550 4256 9555 4312
rect 7852 4254 9555 4256
rect 7852 4252 7858 4254
rect 9489 4251 9555 4254
rect 0 4178 800 4208
rect 2221 4178 2287 4181
rect 3969 4178 4035 4181
rect 4102 4178 4108 4180
rect 0 4176 3802 4178
rect 0 4120 2226 4176
rect 2282 4120 3802 4176
rect 0 4118 3802 4120
rect 0 4088 800 4118
rect 2221 4115 2287 4118
rect 3742 4042 3802 4118
rect 3969 4176 4108 4178
rect 3969 4120 3974 4176
rect 4030 4120 4108 4176
rect 3969 4118 4108 4120
rect 3969 4115 4035 4118
rect 4102 4116 4108 4118
rect 4172 4116 4178 4180
rect 6862 4178 6868 4180
rect 4294 4118 6868 4178
rect 4294 4042 4354 4118
rect 6862 4116 6868 4118
rect 6932 4116 6938 4180
rect 7833 4178 7899 4181
rect 7966 4178 7972 4180
rect 7833 4176 7972 4178
rect 7833 4120 7838 4176
rect 7894 4120 7972 4176
rect 7833 4118 7972 4120
rect 7833 4115 7899 4118
rect 7966 4116 7972 4118
rect 8036 4116 8042 4180
rect 8385 4178 8451 4181
rect 18045 4178 18111 4181
rect 8385 4176 18111 4178
rect 8385 4120 8390 4176
rect 8446 4120 18050 4176
rect 18106 4120 18111 4176
rect 8385 4118 18111 4120
rect 8385 4115 8451 4118
rect 18045 4115 18111 4118
rect 4797 4044 4863 4045
rect 4797 4042 4844 4044
rect 3742 3982 4354 4042
rect 4752 4040 4844 4042
rect 4752 3984 4802 4040
rect 4752 3982 4844 3984
rect 4797 3980 4844 3982
rect 4908 3980 4914 4044
rect 5441 4042 5507 4045
rect 7189 4042 7255 4045
rect 5441 4040 7255 4042
rect 5441 3984 5446 4040
rect 5502 3984 7194 4040
rect 7250 3984 7255 4040
rect 5441 3982 7255 3984
rect 4797 3979 4863 3980
rect 5441 3979 5507 3982
rect 7189 3979 7255 3982
rect 7414 3980 7420 4044
rect 7484 4042 7490 4044
rect 9765 4042 9831 4045
rect 9949 4044 10015 4045
rect 9949 4042 9996 4044
rect 7484 4040 9831 4042
rect 7484 3984 9770 4040
rect 9826 3984 9831 4040
rect 7484 3982 9831 3984
rect 9904 4040 9996 4042
rect 9904 3984 9954 4040
rect 9904 3982 9996 3984
rect 7484 3980 7490 3982
rect 9765 3979 9831 3982
rect 9949 3980 9996 3982
rect 10060 3980 10066 4044
rect 11881 4042 11947 4045
rect 17125 4042 17191 4045
rect 11881 4040 17191 4042
rect 11881 3984 11886 4040
rect 11942 3984 17130 4040
rect 17186 3984 17191 4040
rect 11881 3982 17191 3984
rect 9949 3979 10015 3980
rect 11881 3979 11947 3982
rect 17125 3979 17191 3982
rect 4245 3908 4311 3909
rect 4245 3906 4292 3908
rect 4200 3904 4292 3906
rect 4356 3906 4362 3908
rect 5625 3906 5691 3909
rect 5901 3908 5967 3909
rect 5901 3906 5948 3908
rect 4356 3904 5691 3906
rect 4200 3848 4250 3904
rect 4356 3848 5630 3904
rect 5686 3848 5691 3904
rect 4200 3846 4292 3848
rect 4245 3844 4292 3846
rect 4356 3846 5691 3848
rect 5856 3904 5948 3906
rect 5856 3848 5906 3904
rect 5856 3846 5948 3848
rect 4356 3844 4362 3846
rect 4245 3843 4311 3844
rect 5625 3843 5691 3846
rect 5901 3844 5948 3846
rect 6012 3844 6018 3908
rect 6085 3906 6151 3909
rect 7230 3906 7236 3908
rect 6085 3904 7236 3906
rect 6085 3848 6090 3904
rect 6146 3848 7236 3904
rect 6085 3846 7236 3848
rect 5901 3843 5967 3844
rect 6085 3843 6151 3846
rect 7230 3844 7236 3846
rect 7300 3844 7306 3908
rect 9254 3844 9260 3908
rect 9324 3906 9330 3908
rect 12065 3906 12131 3909
rect 9324 3904 12131 3906
rect 9324 3848 12070 3904
rect 12126 3848 12131 3904
rect 9324 3846 12131 3848
rect 9324 3844 9330 3846
rect 12065 3843 12131 3846
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 933 3770 999 3773
rect 0 3768 999 3770
rect 0 3712 938 3768
rect 994 3712 999 3768
rect 0 3710 999 3712
rect 0 3680 800 3710
rect 933 3707 999 3710
rect 4705 3770 4771 3773
rect 5022 3770 5028 3772
rect 4705 3768 5028 3770
rect 4705 3712 4710 3768
rect 4766 3712 5028 3768
rect 4705 3710 5028 3712
rect 4705 3707 4771 3710
rect 5022 3708 5028 3710
rect 5092 3708 5098 3772
rect 9489 3770 9555 3773
rect 10174 3770 10180 3772
rect 9489 3768 10180 3770
rect 9489 3712 9494 3768
rect 9550 3712 10180 3768
rect 9489 3710 10180 3712
rect 9489 3707 9555 3710
rect 10174 3708 10180 3710
rect 10244 3708 10250 3772
rect 2037 3634 2103 3637
rect 7465 3634 7531 3637
rect 8293 3636 8359 3637
rect 8293 3634 8340 3636
rect 2037 3632 7531 3634
rect 2037 3576 2042 3632
rect 2098 3576 7470 3632
rect 7526 3576 7531 3632
rect 2037 3574 7531 3576
rect 8248 3632 8340 3634
rect 8248 3576 8298 3632
rect 8248 3574 8340 3576
rect 2037 3571 2103 3574
rect 7465 3571 7531 3574
rect 8293 3572 8340 3574
rect 8404 3572 8410 3636
rect 9305 3634 9371 3637
rect 14273 3634 14339 3637
rect 9305 3632 14339 3634
rect 9305 3576 9310 3632
rect 9366 3576 14278 3632
rect 14334 3576 14339 3632
rect 9305 3574 14339 3576
rect 8293 3571 8359 3572
rect 9305 3571 9371 3574
rect 14273 3571 14339 3574
rect 3366 3436 3372 3500
rect 3436 3498 3442 3500
rect 3693 3498 3759 3501
rect 3436 3496 3759 3498
rect 3436 3440 3698 3496
rect 3754 3440 3759 3496
rect 3436 3438 3759 3440
rect 3436 3436 3442 3438
rect 3693 3435 3759 3438
rect 4337 3498 4403 3501
rect 4654 3498 4660 3500
rect 4337 3496 4660 3498
rect 4337 3440 4342 3496
rect 4398 3440 4660 3496
rect 4337 3438 4660 3440
rect 4337 3435 4403 3438
rect 4654 3436 4660 3438
rect 4724 3436 4730 3500
rect 5073 3498 5139 3501
rect 7782 3498 7788 3500
rect 5073 3496 7788 3498
rect 5073 3440 5078 3496
rect 5134 3440 7788 3496
rect 5073 3438 7788 3440
rect 5073 3435 5139 3438
rect 7782 3436 7788 3438
rect 7852 3436 7858 3500
rect 8109 3498 8175 3501
rect 14365 3498 14431 3501
rect 8109 3496 14431 3498
rect 8109 3440 8114 3496
rect 8170 3440 14370 3496
rect 14426 3440 14431 3496
rect 8109 3438 14431 3440
rect 8109 3435 8175 3438
rect 14365 3435 14431 3438
rect 0 3362 800 3392
rect 8661 3362 8727 3365
rect 9029 3362 9095 3365
rect 0 3302 1456 3362
rect 0 3272 800 3302
rect 1396 3090 1456 3302
rect 6686 3302 8586 3362
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 5533 3228 5599 3229
rect 5533 3226 5580 3228
rect 5488 3224 5580 3226
rect 5488 3168 5538 3224
rect 5488 3166 5580 3168
rect 5533 3164 5580 3166
rect 5644 3164 5650 3228
rect 5533 3163 5599 3164
rect 2773 3092 2839 3093
rect 2773 3090 2820 3092
rect 1396 3088 2820 3090
rect 2884 3090 2890 3092
rect 3417 3090 3483 3093
rect 6686 3090 6746 3302
rect 7557 3226 7623 3229
rect 8526 3226 8586 3302
rect 8661 3360 9095 3362
rect 8661 3304 8666 3360
rect 8722 3304 9034 3360
rect 9090 3304 9095 3360
rect 8661 3302 9095 3304
rect 8661 3299 8727 3302
rect 9029 3299 9095 3302
rect 9305 3362 9371 3365
rect 9622 3362 9628 3364
rect 9305 3360 9628 3362
rect 9305 3304 9310 3360
rect 9366 3304 9628 3360
rect 9305 3302 9628 3304
rect 9305 3299 9371 3302
rect 9622 3300 9628 3302
rect 9692 3300 9698 3364
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 9489 3228 9555 3229
rect 9254 3226 9260 3228
rect 7557 3224 8402 3226
rect 7557 3168 7562 3224
rect 7618 3168 8402 3224
rect 7557 3166 8402 3168
rect 8526 3166 9260 3226
rect 7557 3163 7623 3166
rect 8109 3092 8175 3093
rect 8109 3090 8156 3092
rect 1396 3032 2778 3088
rect 1396 3030 2820 3032
rect 2773 3028 2820 3030
rect 2884 3030 2966 3090
rect 3417 3088 6746 3090
rect 3417 3032 3422 3088
rect 3478 3032 6746 3088
rect 3417 3030 6746 3032
rect 8064 3088 8156 3090
rect 8064 3032 8114 3088
rect 8064 3030 8156 3032
rect 2884 3028 2890 3030
rect 2773 3027 2839 3028
rect 3417 3027 3483 3030
rect 8109 3028 8156 3030
rect 8220 3028 8226 3092
rect 8342 3090 8402 3166
rect 9254 3164 9260 3166
rect 9324 3164 9330 3228
rect 9438 3164 9444 3228
rect 9508 3226 9555 3228
rect 9765 3226 9831 3229
rect 9508 3224 9600 3226
rect 9550 3168 9600 3224
rect 9508 3166 9600 3168
rect 9765 3224 10426 3226
rect 9765 3168 9770 3224
rect 9826 3168 10426 3224
rect 9765 3166 10426 3168
rect 9508 3164 9555 3166
rect 9489 3163 9555 3164
rect 9765 3163 9831 3166
rect 10133 3090 10199 3093
rect 8342 3088 10199 3090
rect 8342 3032 10138 3088
rect 10194 3032 10199 3088
rect 8342 3030 10199 3032
rect 10366 3090 10426 3166
rect 17217 3090 17283 3093
rect 10366 3088 17283 3090
rect 10366 3032 17222 3088
rect 17278 3032 17283 3088
rect 10366 3030 17283 3032
rect 8109 3027 8175 3028
rect 10133 3027 10199 3030
rect 17217 3027 17283 3030
rect 0 2954 800 2984
rect 3420 2954 3480 3027
rect 0 2894 3480 2954
rect 5993 2954 6059 2957
rect 13353 2954 13419 2957
rect 5993 2952 13419 2954
rect 5993 2896 5998 2952
rect 6054 2896 13358 2952
rect 13414 2896 13419 2952
rect 5993 2894 13419 2896
rect 0 2864 800 2894
rect 5993 2891 6059 2894
rect 13353 2891 13419 2894
rect 3969 2818 4035 2821
rect 7046 2818 7052 2820
rect 3969 2816 7052 2818
rect 3969 2760 3974 2816
rect 4030 2760 7052 2816
rect 3969 2758 7052 2760
rect 3969 2755 4035 2758
rect 7046 2756 7052 2758
rect 7116 2756 7122 2820
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 2446 2620 2452 2684
rect 2516 2682 2522 2684
rect 6821 2682 6887 2685
rect 7598 2682 7604 2684
rect 2516 2622 3480 2682
rect 2516 2620 2522 2622
rect 0 2546 800 2576
rect 2957 2546 3023 2549
rect 0 2544 3023 2546
rect 0 2488 2962 2544
rect 3018 2488 3023 2544
rect 0 2486 3023 2488
rect 3420 2546 3480 2622
rect 6821 2680 7604 2682
rect 6821 2624 6826 2680
rect 6882 2624 7604 2680
rect 6821 2622 7604 2624
rect 6821 2619 6887 2622
rect 7598 2620 7604 2622
rect 7668 2620 7674 2684
rect 9213 2682 9279 2685
rect 10910 2682 10916 2684
rect 9213 2680 10916 2682
rect 9213 2624 9218 2680
rect 9274 2624 10916 2680
rect 9213 2622 10916 2624
rect 9213 2619 9279 2622
rect 10910 2620 10916 2622
rect 10980 2620 10986 2684
rect 9673 2546 9739 2549
rect 3420 2544 9739 2546
rect 3420 2488 9678 2544
rect 9734 2488 9739 2544
rect 3420 2486 9739 2488
rect 0 2456 800 2486
rect 2957 2483 3023 2486
rect 9673 2483 9739 2486
rect 6729 2410 6795 2413
rect 15929 2410 15995 2413
rect 6729 2408 15995 2410
rect 6729 2352 6734 2408
rect 6790 2352 15934 2408
rect 15990 2352 15995 2408
rect 6729 2350 15995 2352
rect 6729 2347 6795 2350
rect 15929 2347 15995 2350
rect 6637 2274 6703 2277
rect 9806 2274 9812 2276
rect 6637 2272 9812 2274
rect 6637 2216 6642 2272
rect 6698 2216 9812 2272
rect 6637 2214 9812 2216
rect 6637 2211 6703 2214
rect 9806 2212 9812 2214
rect 9876 2212 9882 2276
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 3233 2138 3299 2141
rect 0 2136 3299 2138
rect 0 2080 3238 2136
rect 3294 2080 3299 2136
rect 0 2078 3299 2080
rect 0 2048 800 2078
rect 3233 2075 3299 2078
rect 6678 2076 6684 2140
rect 6748 2138 6754 2140
rect 10961 2138 11027 2141
rect 6748 2136 11027 2138
rect 6748 2080 10966 2136
rect 11022 2080 11027 2136
rect 6748 2078 11027 2080
rect 6748 2076 6754 2078
rect 10961 2075 11027 2078
rect 7966 1940 7972 2004
rect 8036 2002 8042 2004
rect 15193 2002 15259 2005
rect 8036 2000 15259 2002
rect 8036 1944 15198 2000
rect 15254 1944 15259 2000
rect 8036 1942 15259 1944
rect 8036 1940 8042 1942
rect 15193 1939 15259 1942
rect 5901 1866 5967 1869
rect 12065 1866 12131 1869
rect 5901 1864 12131 1866
rect 5901 1808 5906 1864
rect 5962 1808 12070 1864
rect 12126 1808 12131 1864
rect 5901 1806 12131 1808
rect 5901 1803 5967 1806
rect 12065 1803 12131 1806
rect 0 1730 800 1760
rect 4061 1730 4127 1733
rect 0 1728 4127 1730
rect 0 1672 4066 1728
rect 4122 1672 4127 1728
rect 0 1670 4127 1672
rect 0 1640 800 1670
rect 4061 1667 4127 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 9996 14316 10060 14380
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 9444 13908 9508 13972
rect 9812 13832 9876 13836
rect 9812 13776 9826 13832
rect 9826 13776 9876 13832
rect 9812 13772 9876 13776
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 5580 11188 5644 11252
rect 9628 11188 9692 11252
rect 6684 11052 6748 11116
rect 10916 11052 10980 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 3924 9828 3988 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 4476 9692 4540 9756
rect 8156 9692 8220 9756
rect 2820 9556 2884 9620
rect 3372 9420 3436 9484
rect 4660 9420 4724 9484
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 4108 8664 4172 8668
rect 4108 8608 4122 8664
rect 4122 8608 4172 8664
rect 4108 8604 4172 8608
rect 4292 8604 4356 8668
rect 2268 8332 2332 8396
rect 5028 8332 5092 8396
rect 10180 8332 10244 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6868 8120 6932 8124
rect 6868 8064 6882 8120
rect 6882 8064 6932 8120
rect 6868 8060 6932 8064
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 8340 7516 8404 7580
rect 5764 7108 5828 7172
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 2452 6972 2516 7036
rect 4844 6972 4908 7036
rect 7236 6972 7300 7036
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 7420 5884 7484 5948
rect 7052 5748 7116 5812
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 7604 5340 7668 5404
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 5948 4932 6012 4996
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 3924 4660 3988 4724
rect 5764 4524 5828 4588
rect 2268 4388 2332 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 4476 4312 4540 4316
rect 4476 4256 4490 4312
rect 4490 4256 4540 4312
rect 4476 4252 4540 4256
rect 7788 4252 7852 4316
rect 4108 4116 4172 4180
rect 6868 4116 6932 4180
rect 7972 4116 8036 4180
rect 4844 4040 4908 4044
rect 4844 3984 4858 4040
rect 4858 3984 4908 4040
rect 4844 3980 4908 3984
rect 7420 3980 7484 4044
rect 9996 4040 10060 4044
rect 9996 3984 10010 4040
rect 10010 3984 10060 4040
rect 9996 3980 10060 3984
rect 4292 3904 4356 3908
rect 4292 3848 4306 3904
rect 4306 3848 4356 3904
rect 4292 3844 4356 3848
rect 5948 3904 6012 3908
rect 5948 3848 5962 3904
rect 5962 3848 6012 3904
rect 5948 3844 6012 3848
rect 7236 3844 7300 3908
rect 9260 3844 9324 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 5028 3708 5092 3772
rect 10180 3708 10244 3772
rect 8340 3632 8404 3636
rect 8340 3576 8354 3632
rect 8354 3576 8404 3632
rect 8340 3572 8404 3576
rect 3372 3436 3436 3500
rect 4660 3436 4724 3500
rect 7788 3436 7852 3500
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 5580 3224 5644 3228
rect 5580 3168 5594 3224
rect 5594 3168 5644 3224
rect 5580 3164 5644 3168
rect 2820 3088 2884 3092
rect 9628 3300 9692 3364
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 2820 3032 2834 3088
rect 2834 3032 2884 3088
rect 2820 3028 2884 3032
rect 8156 3088 8220 3092
rect 8156 3032 8170 3088
rect 8170 3032 8220 3088
rect 8156 3028 8220 3032
rect 9260 3164 9324 3228
rect 9444 3224 9508 3228
rect 9444 3168 9494 3224
rect 9494 3168 9508 3224
rect 9444 3164 9508 3168
rect 7052 2756 7116 2820
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 2452 2620 2516 2684
rect 7604 2620 7668 2684
rect 10916 2620 10980 2684
rect 9812 2212 9876 2276
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 6684 2076 6748 2140
rect 7972 1940 8036 2004
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 5579 11252 5645 11253
rect 5579 11188 5580 11252
rect 5644 11188 5645 11252
rect 5579 11187 5645 11188
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 2819 9620 2885 9621
rect 2819 9556 2820 9620
rect 2884 9556 2885 9620
rect 2819 9555 2885 9556
rect 2267 8396 2333 8397
rect 2267 8332 2268 8396
rect 2332 8332 2333 8396
rect 2267 8331 2333 8332
rect 2270 4453 2330 8331
rect 2451 7036 2517 7037
rect 2451 6972 2452 7036
rect 2516 6972 2517 7036
rect 2451 6971 2517 6972
rect 2267 4452 2333 4453
rect 2267 4388 2268 4452
rect 2332 4388 2333 4452
rect 2267 4387 2333 4388
rect 2454 2685 2514 6971
rect 2822 3093 2882 9555
rect 3371 9484 3437 9485
rect 3371 9420 3372 9484
rect 3436 9420 3437 9484
rect 3371 9419 3437 9420
rect 3374 3501 3434 9419
rect 3543 9280 3863 10304
rect 3923 9892 3989 9893
rect 3923 9828 3924 9892
rect 3988 9828 3989 9892
rect 3923 9827 3989 9828
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3926 4725 3986 9827
rect 4475 9756 4541 9757
rect 4475 9692 4476 9756
rect 4540 9692 4541 9756
rect 4475 9691 4541 9692
rect 4107 8668 4173 8669
rect 4107 8604 4108 8668
rect 4172 8604 4173 8668
rect 4107 8603 4173 8604
rect 4291 8668 4357 8669
rect 4291 8604 4292 8668
rect 4356 8604 4357 8668
rect 4291 8603 4357 8604
rect 3923 4724 3989 4725
rect 3923 4660 3924 4724
rect 3988 4660 3989 4724
rect 3923 4659 3989 4660
rect 4110 4181 4170 8603
rect 4107 4180 4173 4181
rect 4107 4116 4108 4180
rect 4172 4116 4173 4180
rect 4107 4115 4173 4116
rect 4294 3909 4354 8603
rect 4478 4317 4538 9691
rect 4659 9484 4725 9485
rect 4659 9420 4660 9484
rect 4724 9420 4725 9484
rect 4659 9419 4725 9420
rect 4475 4316 4541 4317
rect 4475 4252 4476 4316
rect 4540 4252 4541 4316
rect 4475 4251 4541 4252
rect 4291 3908 4357 3909
rect 4291 3844 4292 3908
rect 4356 3844 4357 3908
rect 4291 3843 4357 3844
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3371 3500 3437 3501
rect 3371 3436 3372 3500
rect 3436 3436 3437 3500
rect 3371 3435 3437 3436
rect 2819 3092 2885 3093
rect 2819 3028 2820 3092
rect 2884 3028 2885 3092
rect 2819 3027 2885 3028
rect 3543 2752 3863 3776
rect 4662 3501 4722 9419
rect 5027 8396 5093 8397
rect 5027 8332 5028 8396
rect 5092 8332 5093 8396
rect 5027 8331 5093 8332
rect 4843 7036 4909 7037
rect 4843 6972 4844 7036
rect 4908 6972 4909 7036
rect 4843 6971 4909 6972
rect 4846 4045 4906 6971
rect 4843 4044 4909 4045
rect 4843 3980 4844 4044
rect 4908 3980 4909 4044
rect 4843 3979 4909 3980
rect 5030 3773 5090 8331
rect 5027 3772 5093 3773
rect 5027 3708 5028 3772
rect 5092 3708 5093 3772
rect 5027 3707 5093 3708
rect 4659 3500 4725 3501
rect 4659 3436 4660 3500
rect 4724 3436 4725 3500
rect 4659 3435 4725 3436
rect 5582 3229 5642 11187
rect 6142 10912 6462 11936
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 9995 14380 10061 14381
rect 9995 14316 9996 14380
rect 10060 14316 10061 14380
rect 9995 14315 10061 14316
rect 9443 13972 9509 13973
rect 9443 13908 9444 13972
rect 9508 13908 9509 13972
rect 9443 13907 9509 13908
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 6683 11116 6749 11117
rect 6683 11052 6684 11116
rect 6748 11052 6749 11116
rect 6683 11051 6749 11052
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 5763 7172 5829 7173
rect 5763 7108 5764 7172
rect 5828 7108 5829 7172
rect 5763 7107 5829 7108
rect 5766 4589 5826 7107
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 5947 4996 6013 4997
rect 5947 4932 5948 4996
rect 6012 4932 6013 4996
rect 5947 4931 6013 4932
rect 5763 4588 5829 4589
rect 5763 4524 5764 4588
rect 5828 4524 5829 4588
rect 5763 4523 5829 4524
rect 5950 3909 6010 4931
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5947 3908 6013 3909
rect 5947 3844 5948 3908
rect 6012 3844 6013 3908
rect 5947 3843 6013 3844
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5579 3228 5645 3229
rect 5579 3164 5580 3228
rect 5644 3164 5645 3228
rect 5579 3163 5645 3164
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 2451 2684 2517 2685
rect 2451 2620 2452 2684
rect 2516 2620 2517 2684
rect 2451 2619 2517 2620
rect 3543 2128 3863 2688
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 6686 2141 6746 11051
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 6867 8124 6933 8125
rect 6867 8060 6868 8124
rect 6932 8060 6933 8124
rect 6867 8059 6933 8060
rect 6870 4181 6930 8059
rect 7235 7036 7301 7037
rect 7235 6972 7236 7036
rect 7300 6972 7301 7036
rect 7235 6971 7301 6972
rect 7051 5812 7117 5813
rect 7051 5748 7052 5812
rect 7116 5748 7117 5812
rect 7051 5747 7117 5748
rect 6867 4180 6933 4181
rect 6867 4116 6868 4180
rect 6932 4116 6933 4180
rect 6867 4115 6933 4116
rect 7054 2821 7114 5747
rect 7238 3909 7298 6971
rect 7419 5948 7485 5949
rect 7419 5884 7420 5948
rect 7484 5884 7485 5948
rect 7419 5883 7485 5884
rect 7422 4045 7482 5883
rect 7603 5404 7669 5405
rect 7603 5340 7604 5404
rect 7668 5340 7669 5404
rect 7603 5339 7669 5340
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 7235 3908 7301 3909
rect 7235 3844 7236 3908
rect 7300 3844 7301 3908
rect 7235 3843 7301 3844
rect 7051 2820 7117 2821
rect 7051 2756 7052 2820
rect 7116 2756 7117 2820
rect 7051 2755 7117 2756
rect 7606 2685 7666 5339
rect 7787 4316 7853 4317
rect 7787 4252 7788 4316
rect 7852 4252 7853 4316
rect 7787 4251 7853 4252
rect 7790 3501 7850 4251
rect 7971 4180 8037 4181
rect 7971 4116 7972 4180
rect 8036 4116 8037 4180
rect 7971 4115 8037 4116
rect 7787 3500 7853 3501
rect 7787 3436 7788 3500
rect 7852 3436 7853 3500
rect 7787 3435 7853 3436
rect 7603 2684 7669 2685
rect 7603 2620 7604 2684
rect 7668 2620 7669 2684
rect 7603 2619 7669 2620
rect 6683 2140 6749 2141
rect 6683 2076 6684 2140
rect 6748 2076 6749 2140
rect 6683 2075 6749 2076
rect 7974 2005 8034 4115
rect 8158 3093 8218 9691
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8339 7580 8405 7581
rect 8339 7516 8340 7580
rect 8404 7516 8405 7580
rect 8339 7515 8405 7516
rect 8342 3637 8402 7515
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 9259 3908 9325 3909
rect 9259 3844 9260 3908
rect 9324 3844 9325 3908
rect 9259 3843 9325 3844
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8339 3636 8405 3637
rect 8339 3572 8340 3636
rect 8404 3572 8405 3636
rect 8339 3571 8405 3572
rect 8155 3092 8221 3093
rect 8155 3028 8156 3092
rect 8220 3028 8221 3092
rect 8155 3027 8221 3028
rect 8741 2752 9061 3776
rect 9262 3229 9322 3843
rect 9446 3229 9506 13907
rect 9811 13836 9877 13837
rect 9811 13772 9812 13836
rect 9876 13772 9877 13836
rect 9811 13771 9877 13772
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 9630 3365 9690 11187
rect 9627 3364 9693 3365
rect 9627 3300 9628 3364
rect 9692 3300 9693 3364
rect 9627 3299 9693 3300
rect 9259 3228 9325 3229
rect 9259 3164 9260 3228
rect 9324 3164 9325 3228
rect 9259 3163 9325 3164
rect 9443 3228 9509 3229
rect 9443 3164 9444 3228
rect 9508 3164 9509 3228
rect 9443 3163 9509 3164
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 9814 2277 9874 13771
rect 9998 4045 10058 14315
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 10179 8396 10245 8397
rect 10179 8332 10180 8396
rect 10244 8332 10245 8396
rect 10179 8331 10245 8332
rect 9995 4044 10061 4045
rect 9995 3980 9996 4044
rect 10060 3980 10061 4044
rect 9995 3979 10061 3980
rect 10182 3773 10242 8331
rect 10179 3772 10245 3773
rect 10179 3708 10180 3772
rect 10244 3708 10245 3772
rect 10179 3707 10245 3708
rect 10918 2685 10978 11051
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10915 2684 10981 2685
rect 10915 2620 10916 2684
rect 10980 2620 10981 2684
rect 10915 2619 10981 2620
rect 9811 2276 9877 2277
rect 9811 2212 9812 2276
rect 9876 2212 9877 2276
rect 9811 2211 9877 2212
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
rect 7971 2004 8037 2005
rect 7971 1940 7972 2004
rect 8036 1940 8037 2004
rect 7971 1939 8037 1940
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 5888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 17112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 5796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 6716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 8372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 10948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 9108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 6992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 4324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 3220 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19044 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20884 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 1564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3128 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1649977179
transform -1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform -1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform -1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform -1 0 18676 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1649977179
transform -1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1649977179
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_82
timestamp 1649977179
transform 1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1649977179
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1649977179
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_34
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp 1649977179
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1649977179
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_126
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1649977179
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_164
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_213
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_32
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1649977179
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1649977179
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_61
timestamp 1649977179
transform 1 0 6716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1649977179
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1649977179
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_116
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_120
timestamp 1649977179
transform 1 0 12144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1649977179
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_96
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_101
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_107
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1649977179
transform 1 0 13064 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_146
timestamp 1649977179
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_6
timestamp 1649977179
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_10
timestamp 1649977179
transform 1 0 2024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1649977179
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_195
timestamp 1649977179
transform 1 0 19044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1649977179
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1649977179
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp 1649977179
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1649977179
transform 1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_132
timestamp 1649977179
transform 1 0 13248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_166
timestamp 1649977179
transform 1 0 16376 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_170
timestamp 1649977179
transform 1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1649977179
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_35
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1649977179
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1649977179
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_185
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_215
timestamp 1649977179
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1649977179
transform 1 0 7544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1649977179
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_98
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_106
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp 1649977179
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_217
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_6
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp 1649977179
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1649977179
transform 1 0 5520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_63
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1649977179
transform 1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1649977179
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_155
timestamp 1649977179
transform 1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1649977179
transform 1 0 17204 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1649977179
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_16
timestamp 1649977179
transform 1 0 2576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1649977179
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1649977179
transform 1 0 4968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1649977179
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_159
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_213
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_10
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_26
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_99 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1649977179
transform 1 0 19780 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1649977179
transform 1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_200
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_6
timestamp 1649977179
transform 1 0 1656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_23
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_89
timestamp 1649977179
transform 1 0 9292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1649977179
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_153
timestamp 1649977179
transform 1 0 15180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_214
timestamp 1649977179
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_218
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_16
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_20
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_34
timestamp 1649977179
transform 1 0 4232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_99 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_125
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_148
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_213
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_18
timestamp 1649977179
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_72
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_90
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp 1649977179
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1649977179
transform 1 0 14536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_5
timestamp 1649977179
transform 1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1649977179
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_31
timestamp 1649977179
transform 1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_35
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1649977179
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_57
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_61
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_88
timestamp 1649977179
transform 1 0 9200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1649977179
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_6
timestamp 1649977179
transform 1 0 1656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_10
timestamp 1649977179
transform 1 0 2024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_66
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1649977179
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_10
timestamp 1649977179
transform 1 0 2024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_31
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1649977179
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1649977179
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_178
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1649977179
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1649977179
transform 1 0 2208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_24
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_28
timestamp 1649977179
transform 1 0 3680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_32
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_44
timestamp 1649977179
transform 1 0 5152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_61
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_87
timestamp 1649977179
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_141
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1649977179
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_215
timestamp 1649977179
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_5
timestamp 1649977179
transform 1 0 1564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_16
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1649977179
transform 1 0 3036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_42
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_48
timestamp 1649977179
transform 1 0 5520 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_128
timestamp 1649977179
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1649977179
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_38
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_59
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_133
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_145
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1649977179
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_45
timestamp 1649977179
transform 1 0 5244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_98
timestamp 1649977179
transform 1 0 10120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_103
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_112
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 1649977179
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_17
timestamp 1649977179
transform 1 0 2668 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_23
timestamp 1649977179
transform 1 0 3220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_59
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1649977179
transform 1 0 7728 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_77
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_89
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_38
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_47
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_59
timestamp 1649977179
transform 1 0 6532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1649977179
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_75
timestamp 1649977179
transform 1 0 8004 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_87
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_99
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_33
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_49
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_99
timestamp 1649977179
transform 1 0 10212 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_103
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_127
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_17
timestamp 1649977179
transform 1 0 2668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_25
timestamp 1649977179
transform 1 0 3404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_30
timestamp 1649977179
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1649977179
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_70
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_82
timestamp 1649977179
transform 1 0 8648 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_94
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1649977179
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_13
timestamp 1649977179
transform 1 0 2300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_33
timestamp 1649977179
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 1649977179
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_66
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1649977179
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_19
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_31
timestamp 1649977179
transform 1 0 3956 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_40
timestamp 1649977179
transform 1 0 4784 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_52
timestamp 1649977179
transform 1 0 5888 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_64
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1649977179
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_33
timestamp 1649977179
transform 1 0 4140 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_82
timestamp 1649977179
transform 1 0 8648 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_94
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_39
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_47
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_51
timestamp 1649977179
transform 1 0 5796 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_63
timestamp 1649977179
transform 1 0 6900 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_69
timestamp 1649977179
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1649977179
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_23
timestamp 1649977179
transform 1 0 3220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _070_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 2760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 3864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform 1 0 4416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 13156 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 18952 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform -1 0 3404 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform -1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform -1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform -1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1649977179
transform -1 0 3404 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11224 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12696 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21160 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18216 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16100 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15180 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17020 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18400 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20516 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17388 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18492 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15640 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12880 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14812 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13156 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12880 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14076 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12788 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11776 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14260 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21160 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18768 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17112 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_1__127 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3220 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2208 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_1__103
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_1__104
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7452 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4508 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3864 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_7.mux_l2_in_1__105
timestamp 1649977179
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_0__106
timestamp 1649977179
transform -1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_11.mux_l2_in_0__128
timestamp 1649977179
transform -1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_13.mux_l2_in_0__129
timestamp 1649977179
transform 1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6716 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_15.mux_l2_in_0__130
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_0__131
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8096 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_19.mux_l2_in_0__132
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_21.mux_l2_in_0__133
timestamp 1649977179
transform -1 0 9568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_23.mux_l2_in_0__134
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5152 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l1_in_1__135
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5520 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5520 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_27.mux_l2_in_0__136
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9384 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_29.mux_l2_in_0__137
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_1__107
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3312 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_1__118
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform -1 0 2576 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_1__124
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 1932 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2576 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4324 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_7.mux_l2_in_1__125
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l1_in_1__126
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_11.mux_l2_in_0__108
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_13.mux_l2_in_0__109
timestamp 1649977179
transform 1 0 6900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_15.mux_l2_in_0__110
timestamp 1649977179
transform -1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_0__111
timestamp 1649977179
transform -1 0 6716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_19.mux_l2_in_0__112
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_21.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4232 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_23.mux_l2_in_0__114
timestamp 1649977179
transform 1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4876 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_1__115
timestamp 1649977179
transform 1 0 5244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_27.mux_l2_in_0__116
timestamp 1649977179
transform -1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_29.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 8924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_31.mux_l2_in_0__119
timestamp 1649977179
transform -1 0 9568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7452 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_0__120
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_35.mux_l2_in_0__121
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12512 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_37.mux_l2_in_0__122
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_39.mux_l2_in_0__123
timestamp 1649977179
transform 1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
<< labels >>
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 0 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 bottom_right_grid_pin_1_
port 12 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 ccff_head
port 13 nsew signal input
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 ccff_tail
port 14 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 15 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 16 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 17 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 18 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 19 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 20 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 21 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 22 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 23 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 24 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 25 nsew signal input
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 26 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 27 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 28 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 29 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 30 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 31 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 32 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 33 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 34 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 35 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 36 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 37 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 38 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 39 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 40 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 41 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 42 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 43 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 44 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 45 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 46 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 47 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 48 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 49 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 50 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 51 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 52 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 53 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 54 nsew signal tristate
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 55 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 56 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 57 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 58 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 59 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 60 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 61 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 62 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 63 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 64 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 65 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 66 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 67 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 68 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 69 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 70 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 71 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 72 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 73 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 74 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 75 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 76 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 77 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 78 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 79 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 80 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 81 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 82 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 83 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 84 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 85 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 86 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 87 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 88 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 89 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 90 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 91 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 92 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 93 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 94 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 95 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 96 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 97 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 98 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 99 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 100 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 101 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 102 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 left_top_grid_pin_1_
port 103 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 104 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
