magic
tech sky130A
magscale 1 2
timestamp 1681041352
<< viali >>
rect 13829 54281 13863 54315
rect 18981 54281 19015 54315
rect 2421 54213 2455 54247
rect 5089 54213 5123 54247
rect 3433 54145 3467 54179
rect 6009 54145 6043 54179
rect 8401 54145 8435 54179
rect 9597 54145 9631 54179
rect 12173 54145 12207 54179
rect 14473 54145 14507 54179
rect 15117 54145 15151 54179
rect 15393 54145 15427 54179
rect 17049 54145 17083 54179
rect 17325 54145 17359 54179
rect 17877 54145 17911 54179
rect 18153 54145 18187 54179
rect 19441 54145 19475 54179
rect 21005 54145 21039 54179
rect 21281 54145 21315 54179
rect 22293 54145 22327 54179
rect 22569 54145 22603 54179
rect 24041 54145 24075 54179
rect 24685 54145 24719 54179
rect 25329 54145 25363 54179
rect 7849 54077 7883 54111
rect 9873 54077 9907 54111
rect 12633 54077 12667 54111
rect 19717 54077 19751 54111
rect 23121 54077 23155 54111
rect 14933 54009 14967 54043
rect 20821 54009 20855 54043
rect 14289 53941 14323 53975
rect 16865 53941 16899 53975
rect 17693 53941 17727 53975
rect 22109 53941 22143 53975
rect 23397 53941 23431 53975
rect 1777 53601 1811 53635
rect 4169 53601 4203 53635
rect 6929 53601 6963 53635
rect 11253 53601 11287 53635
rect 2973 53533 3007 53567
rect 5365 53533 5399 53567
rect 8033 53533 8067 53567
rect 10793 53533 10827 53567
rect 22569 53533 22603 53567
rect 23213 53533 23247 53567
rect 23765 53533 23799 53567
rect 24685 53533 24719 53567
rect 23029 53465 23063 53499
rect 22385 53397 22419 53431
rect 23949 53397 23983 53431
rect 25329 53397 25363 53431
rect 5181 53193 5215 53227
rect 22661 53193 22695 53227
rect 23305 53193 23339 53227
rect 23397 53193 23431 53227
rect 25053 53193 25087 53227
rect 25329 53193 25363 53227
rect 5365 53057 5399 53091
rect 24041 53057 24075 53091
rect 24777 53057 24811 53091
rect 25513 52921 25547 52955
rect 23857 52853 23891 52887
rect 24593 52853 24627 52887
rect 6561 52649 6595 52683
rect 24501 52649 24535 52683
rect 23857 52581 23891 52615
rect 24961 52513 24995 52547
rect 6745 52445 6779 52479
rect 24041 52445 24075 52479
rect 25237 52377 25271 52411
rect 24133 52105 24167 52139
rect 24593 51969 24627 52003
rect 25329 51969 25363 52003
rect 24409 51765 24443 51799
rect 25145 51765 25179 51799
rect 8309 51561 8343 51595
rect 9229 51561 9263 51595
rect 7573 51493 7607 51527
rect 8493 51357 8527 51391
rect 9413 51357 9447 51391
rect 7757 51289 7791 51323
rect 24593 51289 24627 51323
rect 25237 51289 25271 51323
rect 25145 51221 25179 51255
rect 24593 50881 24627 50915
rect 25237 50881 25271 50915
rect 25145 50677 25179 50711
rect 7757 50473 7791 50507
rect 8401 50473 8435 50507
rect 9597 50473 9631 50507
rect 7573 50405 7607 50439
rect 8033 50269 8067 50303
rect 9505 50269 9539 50303
rect 25421 50133 25455 50167
rect 25053 49725 25087 49759
rect 25329 49725 25363 49759
rect 10701 49317 10735 49351
rect 11713 49317 11747 49351
rect 10517 49113 10551 49147
rect 11529 49113 11563 49147
rect 24777 49113 24811 49147
rect 25237 49113 25271 49147
rect 25145 49045 25179 49079
rect 6653 48841 6687 48875
rect 8125 48637 8159 48671
rect 8401 48637 8435 48671
rect 8677 48501 8711 48535
rect 8953 48501 8987 48535
rect 25421 48501 25455 48535
rect 10368 48093 10402 48127
rect 24041 48093 24075 48127
rect 25237 48093 25271 48127
rect 10471 47957 10505 47991
rect 23397 47957 23431 47991
rect 25145 47957 25179 47991
rect 9873 47753 9907 47787
rect 10149 47685 10183 47719
rect 9413 47617 9447 47651
rect 24869 47617 24903 47651
rect 25329 47617 25363 47651
rect 9505 47413 9539 47447
rect 25145 47413 25179 47447
rect 11656 47005 11690 47039
rect 11759 46937 11793 46971
rect 25421 46869 25455 46903
rect 10333 46665 10367 46699
rect 11069 46665 11103 46699
rect 14105 46597 14139 46631
rect 10793 46529 10827 46563
rect 12576 46529 12610 46563
rect 13921 46529 13955 46563
rect 25329 46529 25363 46563
rect 15761 46461 15795 46495
rect 10609 46325 10643 46359
rect 12679 46325 12713 46359
rect 25145 46325 25179 46359
rect 7941 46121 7975 46155
rect 8401 45985 8435 46019
rect 16221 45985 16255 46019
rect 16681 45985 16715 46019
rect 8585 45917 8619 45951
rect 13312 45917 13346 45951
rect 24869 45917 24903 45951
rect 25329 45917 25363 45951
rect 16497 45849 16531 45883
rect 13415 45781 13449 45815
rect 25145 45781 25179 45815
rect 12909 45509 12943 45543
rect 12725 45441 12759 45475
rect 14565 45373 14599 45407
rect 25421 45237 25455 45271
rect 9137 45033 9171 45067
rect 17049 44897 17083 44931
rect 17509 44897 17543 44931
rect 10885 44829 10919 44863
rect 25329 44829 25363 44863
rect 10609 44761 10643 44795
rect 17325 44761 17359 44795
rect 11161 44693 11195 44727
rect 11345 44693 11379 44727
rect 25145 44693 25179 44727
rect 9597 44489 9631 44523
rect 9137 44353 9171 44387
rect 11069 44353 11103 44387
rect 11529 44353 11563 44387
rect 24777 44353 24811 44387
rect 25237 44353 25271 44387
rect 8953 44285 8987 44319
rect 10609 44149 10643 44183
rect 10977 44149 11011 44183
rect 25145 44149 25179 44183
rect 21833 43809 21867 43843
rect 22109 43741 22143 43775
rect 20361 43605 20395 43639
rect 22385 43605 22419 43639
rect 25421 43605 25455 43639
rect 25237 43265 25271 43299
rect 25053 43129 25087 43163
rect 9781 42721 9815 42755
rect 10241 42721 10275 42755
rect 9597 42653 9631 42687
rect 24777 42585 24811 42619
rect 25237 42585 25271 42619
rect 25145 42517 25179 42551
rect 9413 42313 9447 42347
rect 10885 42245 10919 42279
rect 11161 42109 11195 42143
rect 11529 41973 11563 42007
rect 11713 41973 11747 42007
rect 25421 41973 25455 42007
rect 10885 41769 10919 41803
rect 10425 41633 10459 41667
rect 10241 41565 10275 41599
rect 25237 41565 25271 41599
rect 25053 41497 25087 41531
rect 24869 41089 24903 41123
rect 25329 41089 25363 41123
rect 25145 40885 25179 40919
rect 25513 40341 25547 40375
rect 25145 40137 25179 40171
rect 25329 40001 25363 40035
rect 24869 39389 24903 39423
rect 25329 39389 25363 39423
rect 25145 39253 25179 39287
rect 25421 38709 25455 38743
rect 25329 38301 25363 38335
rect 25145 38165 25179 38199
rect 8677 37961 8711 37995
rect 8861 37825 8895 37859
rect 24777 37825 24811 37859
rect 25237 37825 25271 37859
rect 25145 37621 25179 37655
rect 25421 37077 25455 37111
rect 25237 36737 25271 36771
rect 25145 36533 25179 36567
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 25145 35989 25179 36023
rect 22477 35785 22511 35819
rect 11529 35717 11563 35751
rect 21189 35717 21223 35751
rect 9413 35649 9447 35683
rect 20453 35649 20487 35683
rect 21097 35649 21131 35683
rect 22385 35649 22419 35683
rect 9689 35581 9723 35615
rect 11161 35581 11195 35615
rect 21281 35581 21315 35615
rect 22569 35581 22603 35615
rect 22017 35513 22051 35547
rect 11805 35445 11839 35479
rect 20729 35445 20763 35479
rect 25421 35445 25455 35479
rect 21833 35241 21867 35275
rect 23305 35105 23339 35139
rect 23213 35037 23247 35071
rect 25329 35037 25363 35071
rect 22385 34969 22419 35003
rect 23121 34969 23155 35003
rect 22753 34901 22787 34935
rect 25145 34901 25179 34935
rect 25145 34697 25179 34731
rect 24869 34561 24903 34595
rect 25329 34561 25363 34595
rect 21373 34357 21407 34391
rect 9137 34153 9171 34187
rect 21649 34153 21683 34187
rect 14749 34017 14783 34051
rect 23121 34017 23155 34051
rect 23397 34017 23431 34051
rect 9321 33949 9355 33983
rect 19441 33949 19475 33983
rect 24869 33949 24903 33983
rect 25329 33949 25363 33983
rect 15577 33881 15611 33915
rect 15853 33881 15887 33915
rect 19717 33881 19751 33915
rect 21189 33813 21223 33847
rect 23765 33813 23799 33847
rect 25145 33813 25179 33847
rect 21649 33609 21683 33643
rect 23765 33609 23799 33643
rect 22293 33541 22327 33575
rect 25329 33473 25363 33507
rect 21005 33405 21039 33439
rect 21281 33405 21315 33439
rect 22017 33405 22051 33439
rect 19533 33269 19567 33303
rect 24225 33269 24259 33303
rect 24317 33269 24351 33303
rect 24593 33269 24627 33303
rect 24869 33269 24903 33303
rect 25145 33269 25179 33303
rect 16773 33065 16807 33099
rect 22293 33065 22327 33099
rect 17049 32997 17083 33031
rect 16221 32929 16255 32963
rect 16589 32929 16623 32963
rect 24041 32929 24075 32963
rect 24777 32929 24811 32963
rect 16037 32861 16071 32895
rect 24869 32861 24903 32895
rect 15945 32793 15979 32827
rect 19901 32793 19935 32827
rect 20729 32793 20763 32827
rect 23765 32793 23799 32827
rect 15577 32725 15611 32759
rect 19625 32725 19659 32759
rect 24961 32725 24995 32759
rect 25329 32725 25363 32759
rect 16865 32521 16899 32555
rect 16313 32453 16347 32487
rect 20545 32453 20579 32487
rect 22109 32385 22143 32419
rect 22937 32385 22971 32419
rect 23489 32385 23523 32419
rect 15485 32317 15519 32351
rect 20821 32317 20855 32351
rect 23765 32317 23799 32351
rect 17049 32181 17083 32215
rect 19073 32181 19107 32215
rect 21097 32181 21131 32215
rect 21649 32181 21683 32215
rect 25237 32181 25271 32215
rect 15577 31909 15611 31943
rect 23029 31909 23063 31943
rect 25145 31909 25179 31943
rect 16037 31841 16071 31875
rect 16221 31841 16255 31875
rect 18521 31841 18555 31875
rect 19717 31841 19751 31875
rect 21189 31841 21223 31875
rect 22109 31841 22143 31875
rect 22201 31841 22235 31875
rect 23489 31841 23523 31875
rect 23581 31841 23615 31875
rect 16773 31773 16807 31807
rect 19441 31773 19475 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 17049 31705 17083 31739
rect 15945 31637 15979 31671
rect 18797 31637 18831 31671
rect 21649 31637 21683 31671
rect 22017 31637 22051 31671
rect 22661 31637 22695 31671
rect 23397 31637 23431 31671
rect 24041 31637 24075 31671
rect 15577 31433 15611 31467
rect 16405 31433 16439 31467
rect 19165 31433 19199 31467
rect 20545 31433 20579 31467
rect 14933 31365 14967 31399
rect 21281 31365 21315 31399
rect 21557 31365 21591 31399
rect 22753 31365 22787 31399
rect 17417 31297 17451 31331
rect 19809 31297 19843 31331
rect 20453 31297 20487 31331
rect 22477 31297 22511 31331
rect 25329 31297 25363 31331
rect 15209 31229 15243 31263
rect 17693 31229 17727 31263
rect 20637 31229 20671 31263
rect 20085 31161 20119 31195
rect 13461 31093 13495 31127
rect 15761 31093 15795 31127
rect 16773 31093 16807 31127
rect 19441 31093 19475 31127
rect 24225 31093 24259 31127
rect 24593 31093 24627 31127
rect 25145 31093 25179 31127
rect 9321 30889 9355 30923
rect 15669 30889 15703 30923
rect 15853 30889 15887 30923
rect 16773 30889 16807 30923
rect 22477 30889 22511 30923
rect 25513 30889 25547 30923
rect 18521 30753 18555 30787
rect 20729 30753 20763 30787
rect 9137 30685 9171 30719
rect 15301 30685 15335 30719
rect 14565 30617 14599 30651
rect 18245 30617 18279 30651
rect 21005 30617 21039 30651
rect 24593 30617 24627 30651
rect 18797 30549 18831 30583
rect 20269 30549 20303 30583
rect 22845 30549 22879 30583
rect 23213 30549 23247 30583
rect 20269 30345 20303 30379
rect 15025 30277 15059 30311
rect 20361 30277 20395 30311
rect 22477 30277 22511 30311
rect 8953 30209 8987 30243
rect 13553 30209 13587 30243
rect 15853 30209 15887 30243
rect 21465 30209 21499 30243
rect 22385 30209 22419 30243
rect 13277 30141 13311 30175
rect 14197 30141 14231 30175
rect 15577 30141 15611 30175
rect 15761 30141 15795 30175
rect 16773 30141 16807 30175
rect 20453 30141 20487 30175
rect 22569 30141 22603 30175
rect 23305 30141 23339 30175
rect 23581 30141 23615 30175
rect 25053 30141 25087 30175
rect 9137 30073 9171 30107
rect 11805 30005 11839 30039
rect 16221 30005 16255 30039
rect 16957 30005 16991 30039
rect 18889 30005 18923 30039
rect 19901 30005 19935 30039
rect 22017 30005 22051 30039
rect 12909 29801 12943 29835
rect 13461 29801 13495 29835
rect 16313 29801 16347 29835
rect 24593 29801 24627 29835
rect 20177 29733 20211 29767
rect 25145 29733 25179 29767
rect 11161 29665 11195 29699
rect 15301 29665 15335 29699
rect 15485 29665 15519 29699
rect 16497 29665 16531 29699
rect 20637 29665 20671 29699
rect 20729 29665 20763 29699
rect 15577 29597 15611 29631
rect 18797 29597 18831 29631
rect 23397 29597 23431 29631
rect 23857 29597 23891 29631
rect 25329 29597 25363 29631
rect 11437 29529 11471 29563
rect 18521 29529 18555 29563
rect 22937 29529 22971 29563
rect 13185 29461 13219 29495
rect 13645 29461 13679 29495
rect 15945 29461 15979 29495
rect 17049 29461 17083 29495
rect 19441 29461 19475 29495
rect 20545 29461 20579 29495
rect 23213 29461 23247 29495
rect 24041 29461 24075 29495
rect 24501 29461 24535 29495
rect 9505 29257 9539 29291
rect 12541 29257 12575 29291
rect 12633 29257 12667 29291
rect 15117 29257 15151 29291
rect 15945 29257 15979 29291
rect 16037 29257 16071 29291
rect 17325 29257 17359 29291
rect 17877 29257 17911 29291
rect 19165 29257 19199 29291
rect 19257 29257 19291 29291
rect 23949 29257 23983 29291
rect 25421 29257 25455 29291
rect 9965 29189 9999 29223
rect 19993 29189 20027 29223
rect 9873 29121 9907 29155
rect 13369 29121 13403 29155
rect 17233 29121 17267 29155
rect 21833 29121 21867 29155
rect 22201 29121 22235 29155
rect 24041 29121 24075 29155
rect 25329 29121 25363 29155
rect 10057 29053 10091 29087
rect 12817 29053 12851 29087
rect 16129 29053 16163 29087
rect 17417 29053 17451 29087
rect 19349 29053 19383 29087
rect 23029 29053 23063 29087
rect 24133 29053 24167 29087
rect 24961 29053 24995 29087
rect 12173 28985 12207 29019
rect 15577 28985 15611 29019
rect 16865 28985 16899 29019
rect 18061 28985 18095 29019
rect 18797 28985 18831 29019
rect 23581 28985 23615 29019
rect 13626 28917 13660 28951
rect 9137 28713 9171 28747
rect 18889 28713 18923 28747
rect 22385 28713 22419 28747
rect 22845 28645 22879 28679
rect 15393 28577 15427 28611
rect 15853 28577 15887 28611
rect 17417 28577 17451 28611
rect 20085 28577 20119 28611
rect 23397 28577 23431 28611
rect 25145 28577 25179 28611
rect 10885 28509 10919 28543
rect 11437 28509 11471 28543
rect 17141 28509 17175 28543
rect 20637 28509 20671 28543
rect 24961 28509 24995 28543
rect 25053 28509 25087 28543
rect 10609 28441 10643 28475
rect 11713 28441 11747 28475
rect 15301 28441 15335 28475
rect 20913 28441 20947 28475
rect 23305 28441 23339 28475
rect 13185 28373 13219 28407
rect 13553 28373 13587 28407
rect 14841 28373 14875 28407
rect 15209 28373 15243 28407
rect 16129 28373 16163 28407
rect 16313 28373 16347 28407
rect 19441 28373 19475 28407
rect 19809 28373 19843 28407
rect 19901 28373 19935 28407
rect 23213 28373 23247 28407
rect 23949 28373 23983 28407
rect 24133 28373 24167 28407
rect 24593 28373 24627 28407
rect 13737 28169 13771 28203
rect 15577 28169 15611 28203
rect 16497 28169 16531 28203
rect 19901 28169 19935 28203
rect 22477 28169 22511 28203
rect 11069 28101 11103 28135
rect 17233 28101 17267 28135
rect 22385 28101 22419 28135
rect 25237 28101 25271 28135
rect 15669 28033 15703 28067
rect 16313 28033 16347 28067
rect 17325 28033 17359 28067
rect 21281 28033 21315 28067
rect 11713 27965 11747 27999
rect 11989 27965 12023 27999
rect 15761 27965 15795 27999
rect 17417 27965 17451 27999
rect 18061 27965 18095 27999
rect 18981 27965 19015 27999
rect 20453 27965 20487 27999
rect 22569 27965 22603 27999
rect 24685 27965 24719 27999
rect 24961 27965 24995 27999
rect 19349 27897 19383 27931
rect 13461 27829 13495 27863
rect 15209 27829 15243 27863
rect 16865 27829 16899 27863
rect 18521 27829 18555 27863
rect 18705 27829 18739 27863
rect 21557 27829 21591 27863
rect 22017 27829 22051 27863
rect 23213 27829 23247 27863
rect 25421 27829 25455 27863
rect 12007 27625 12041 27659
rect 21391 27625 21425 27659
rect 22109 27625 22143 27659
rect 23593 27625 23627 27659
rect 12265 27489 12299 27523
rect 13553 27489 13587 27523
rect 15853 27489 15887 27523
rect 18061 27489 18095 27523
rect 21649 27489 21683 27523
rect 23857 27489 23891 27523
rect 25053 27489 25087 27523
rect 25145 27489 25179 27523
rect 12633 27421 12667 27455
rect 13461 27421 13495 27455
rect 17877 27421 17911 27455
rect 24225 27421 24259 27455
rect 24961 27421 24995 27455
rect 13369 27353 13403 27387
rect 15669 27353 15703 27387
rect 10517 27285 10551 27319
rect 13001 27285 13035 27319
rect 15209 27285 15243 27319
rect 15577 27285 15611 27319
rect 16221 27285 16255 27319
rect 16405 27285 16439 27319
rect 17509 27285 17543 27319
rect 17969 27285 18003 27319
rect 19901 27285 19935 27319
rect 24593 27285 24627 27319
rect 11069 27081 11103 27115
rect 15669 27081 15703 27115
rect 22753 27081 22787 27115
rect 22845 27081 22879 27115
rect 25329 27081 25363 27115
rect 14565 27013 14599 27047
rect 15761 27013 15795 27047
rect 19441 27013 19475 27047
rect 9321 26945 9355 26979
rect 14841 26945 14875 26979
rect 9597 26877 9631 26911
rect 15853 26877 15887 26911
rect 19717 26877 19751 26911
rect 23029 26877 23063 26911
rect 23581 26877 23615 26911
rect 23857 26877 23891 26911
rect 22385 26809 22419 26843
rect 11529 26741 11563 26775
rect 13093 26741 13127 26775
rect 15301 26741 15335 26775
rect 17969 26741 18003 26775
rect 20085 26741 20119 26775
rect 21833 26741 21867 26775
rect 22017 26741 22051 26775
rect 10885 26537 10919 26571
rect 15669 26537 15703 26571
rect 17233 26537 17267 26571
rect 21189 26537 21223 26571
rect 24041 26537 24075 26571
rect 11345 26469 11379 26503
rect 14289 26469 14323 26503
rect 17049 26469 17083 26503
rect 21465 26469 21499 26503
rect 22661 26469 22695 26503
rect 24593 26469 24627 26503
rect 9137 26401 9171 26435
rect 14841 26401 14875 26435
rect 15393 26401 15427 26435
rect 16129 26401 16163 26435
rect 16221 26401 16255 26435
rect 16773 26401 16807 26435
rect 16957 26401 16991 26435
rect 19717 26401 19751 26435
rect 23213 26401 23247 26435
rect 25145 26401 25179 26435
rect 19441 26333 19475 26367
rect 23121 26333 23155 26367
rect 23857 26333 23891 26367
rect 9413 26265 9447 26299
rect 11253 26265 11287 26299
rect 14657 26265 14691 26299
rect 16037 26265 16071 26299
rect 22385 26265 22419 26299
rect 23029 26265 23063 26299
rect 25053 26265 25087 26299
rect 14749 26197 14783 26231
rect 18245 26197 18279 26231
rect 24961 26197 24995 26231
rect 12449 25993 12483 26027
rect 12909 25993 12943 26027
rect 18153 25993 18187 26027
rect 22477 25993 22511 26027
rect 13921 25925 13955 25959
rect 15301 25925 15335 25959
rect 18245 25925 18279 25959
rect 22385 25925 22419 25959
rect 12541 25857 12575 25891
rect 13829 25857 13863 25891
rect 15209 25857 15243 25891
rect 16037 25857 16071 25891
rect 16865 25857 16899 25891
rect 23489 25857 23523 25891
rect 23949 25857 23983 25891
rect 12265 25789 12299 25823
rect 13645 25789 13679 25823
rect 15393 25789 15427 25823
rect 17417 25789 17451 25823
rect 18429 25789 18463 25823
rect 22569 25789 22603 25823
rect 25145 25789 25179 25823
rect 14289 25721 14323 25755
rect 14841 25653 14875 25687
rect 17049 25653 17083 25687
rect 17785 25653 17819 25687
rect 19073 25653 19107 25687
rect 21557 25653 21591 25687
rect 22017 25653 22051 25687
rect 23305 25653 23339 25687
rect 14289 25449 14323 25483
rect 17141 25449 17175 25483
rect 21741 25449 21775 25483
rect 24501 25449 24535 25483
rect 18153 25381 18187 25415
rect 19349 25381 19383 25415
rect 20361 25381 20395 25415
rect 21005 25381 21039 25415
rect 24593 25381 24627 25415
rect 25145 25381 25179 25415
rect 14841 25313 14875 25347
rect 16313 25313 16347 25347
rect 12633 25245 12667 25279
rect 16957 25245 16991 25279
rect 17601 25245 17635 25279
rect 19901 25245 19935 25279
rect 20821 25245 20855 25279
rect 21557 25245 21591 25279
rect 22661 25245 22695 25279
rect 25329 25245 25363 25279
rect 12357 25177 12391 25211
rect 16129 25177 16163 25211
rect 19717 25177 19751 25211
rect 23857 25177 23891 25211
rect 10885 25109 10919 25143
rect 13001 25109 13035 25143
rect 14657 25109 14691 25143
rect 14749 25109 14783 25143
rect 15301 25109 15335 25143
rect 15761 25109 15795 25143
rect 16221 25109 16255 25143
rect 17785 25109 17819 25143
rect 18337 25109 18371 25143
rect 18705 25109 18739 25143
rect 24869 25109 24903 25143
rect 17233 24905 17267 24939
rect 18429 24905 18463 24939
rect 12081 24837 12115 24871
rect 22477 24837 22511 24871
rect 11989 24769 12023 24803
rect 14749 24769 14783 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 17325 24769 17359 24803
rect 18521 24769 18555 24803
rect 19073 24769 19107 24803
rect 22569 24769 22603 24803
rect 10885 24701 10919 24735
rect 11161 24701 11195 24735
rect 11897 24701 11931 24735
rect 13001 24701 13035 24735
rect 14473 24701 14507 24735
rect 17417 24701 17451 24735
rect 18613 24701 18647 24735
rect 19717 24701 19751 24735
rect 19993 24701 20027 24735
rect 21465 24701 21499 24735
rect 22753 24701 22787 24735
rect 23581 24701 23615 24735
rect 23857 24701 23891 24735
rect 25329 24701 25363 24735
rect 12449 24633 12483 24667
rect 16865 24633 16899 24667
rect 23213 24633 23247 24667
rect 9413 24565 9447 24599
rect 15485 24565 15519 24599
rect 18061 24565 18095 24599
rect 19349 24565 19383 24599
rect 22109 24565 22143 24599
rect 13737 24361 13771 24395
rect 24041 24361 24075 24395
rect 25421 24361 25455 24395
rect 18153 24293 18187 24327
rect 11989 24225 12023 24259
rect 14105 24225 14139 24259
rect 18705 24225 18739 24259
rect 21189 24225 21223 24259
rect 21925 24225 21959 24259
rect 24593 24225 24627 24259
rect 9137 24157 9171 24191
rect 18521 24157 18555 24191
rect 18613 24157 18647 24191
rect 9413 24089 9447 24123
rect 11253 24089 11287 24123
rect 11437 24089 11471 24123
rect 12265 24089 12299 24123
rect 17693 24089 17727 24123
rect 20913 24089 20947 24123
rect 22201 24089 22235 24123
rect 10885 24021 10919 24055
rect 16405 24021 16439 24055
rect 19441 24021 19475 24055
rect 21557 24021 21591 24055
rect 23673 24021 23707 24055
rect 10057 23817 10091 23851
rect 10425 23817 10459 23851
rect 14749 23817 14783 23851
rect 17233 23817 17267 23851
rect 17325 23817 17359 23851
rect 18705 23817 18739 23851
rect 19993 23817 20027 23851
rect 20913 23817 20947 23851
rect 22937 23817 22971 23851
rect 24961 23817 24995 23851
rect 13645 23749 13679 23783
rect 14841 23749 14875 23783
rect 18521 23749 18555 23783
rect 21557 23749 21591 23783
rect 10793 23681 10827 23715
rect 18061 23681 18095 23715
rect 19625 23681 19659 23715
rect 20821 23681 20855 23715
rect 22201 23681 22235 23715
rect 8033 23613 8067 23647
rect 8309 23613 8343 23647
rect 10885 23613 10919 23647
rect 10977 23613 11011 23647
rect 13737 23613 13771 23647
rect 13829 23613 13863 23647
rect 14565 23613 14599 23647
rect 15669 23613 15703 23647
rect 17417 23613 17451 23647
rect 19441 23613 19475 23647
rect 19533 23613 19567 23647
rect 21005 23613 21039 23647
rect 23213 23613 23247 23647
rect 23489 23613 23523 23647
rect 9781 23545 9815 23579
rect 15209 23545 15243 23579
rect 18245 23545 18279 23579
rect 20453 23545 20487 23579
rect 22385 23545 22419 23579
rect 13277 23477 13311 23511
rect 16865 23477 16899 23511
rect 18981 23477 19015 23511
rect 25237 23477 25271 23511
rect 9137 23273 9171 23307
rect 10241 23273 10275 23307
rect 14381 23273 14415 23307
rect 15853 23273 15887 23307
rect 18613 23205 18647 23239
rect 9689 23137 9723 23171
rect 11713 23137 11747 23171
rect 11805 23137 11839 23171
rect 13553 23137 13587 23171
rect 15301 23137 15335 23171
rect 18061 23137 18095 23171
rect 18981 23137 19015 23171
rect 20085 23137 20119 23171
rect 20913 23137 20947 23171
rect 23397 23137 23431 23171
rect 25145 23137 25179 23171
rect 11621 23069 11655 23103
rect 13461 23069 13495 23103
rect 14197 23069 14231 23103
rect 15117 23069 15151 23103
rect 18153 23069 18187 23103
rect 18245 23069 18279 23103
rect 19901 23069 19935 23103
rect 21649 23069 21683 23103
rect 23857 23069 23891 23103
rect 25053 23069 25087 23103
rect 9505 23001 9539 23035
rect 15209 23001 15243 23035
rect 24961 23001 24995 23035
rect 9597 22933 9631 22967
rect 11253 22933 11287 22967
rect 13001 22933 13035 22967
rect 13369 22933 13403 22967
rect 14749 22933 14783 22967
rect 19533 22933 19567 22967
rect 19993 22933 20027 22967
rect 21833 22933 21867 22967
rect 24593 22933 24627 22967
rect 8125 22729 8159 22763
rect 14473 22729 14507 22763
rect 17049 22729 17083 22763
rect 18705 22729 18739 22763
rect 19717 22729 19751 22763
rect 21189 22729 21223 22763
rect 9597 22661 9631 22695
rect 12633 22661 12667 22695
rect 14565 22661 14599 22695
rect 9873 22593 9907 22627
rect 12357 22593 12391 22627
rect 16865 22593 16899 22627
rect 18889 22593 18923 22627
rect 21097 22593 21131 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 10149 22525 10183 22559
rect 21281 22525 21315 22559
rect 22845 22525 22879 22559
rect 24777 22525 24811 22559
rect 14105 22389 14139 22423
rect 20453 22389 20487 22423
rect 20729 22389 20763 22423
rect 23765 22185 23799 22219
rect 10885 22049 10919 22083
rect 12081 22049 12115 22083
rect 12265 22049 12299 22083
rect 14933 22049 14967 22083
rect 15117 22049 15151 22083
rect 16129 22049 16163 22083
rect 19901 22049 19935 22083
rect 21097 22049 21131 22083
rect 25145 22049 25179 22083
rect 23305 21981 23339 22015
rect 23949 21981 23983 22015
rect 24961 21981 24995 22015
rect 25053 21981 25087 22015
rect 12357 21913 12391 21947
rect 16405 21913 16439 21947
rect 18245 21913 18279 21947
rect 23029 21913 23063 21947
rect 8953 21845 8987 21879
rect 10425 21845 10459 21879
rect 10977 21845 11011 21879
rect 11069 21845 11103 21879
rect 11437 21845 11471 21879
rect 12725 21845 12759 21879
rect 15209 21845 15243 21879
rect 15577 21845 15611 21879
rect 17877 21845 17911 21879
rect 19993 21845 20027 21879
rect 20085 21845 20119 21879
rect 20453 21845 20487 21879
rect 21557 21845 21591 21879
rect 24593 21845 24627 21879
rect 8677 21641 8711 21675
rect 9965 21641 9999 21675
rect 10425 21641 10459 21675
rect 11713 21641 11747 21675
rect 19809 21641 19843 21675
rect 21189 21641 21223 21675
rect 22477 21641 22511 21675
rect 10885 21573 10919 21607
rect 15761 21573 15795 21607
rect 21373 21573 21407 21607
rect 9505 21505 9539 21539
rect 9597 21505 9631 21539
rect 10793 21505 10827 21539
rect 14841 21505 14875 21539
rect 18705 21505 18739 21539
rect 19901 21505 19935 21539
rect 20729 21505 20763 21539
rect 22385 21505 22419 21539
rect 25053 21505 25087 21539
rect 6929 21437 6963 21471
rect 7205 21437 7239 21471
rect 9321 21437 9355 21471
rect 10977 21437 11011 21471
rect 14565 21437 14599 21471
rect 19717 21437 19751 21471
rect 22661 21437 22695 21471
rect 24777 21437 24811 21471
rect 15577 21369 15611 21403
rect 18889 21369 18923 21403
rect 13093 21301 13127 21335
rect 15117 21301 15151 21335
rect 19165 21301 19199 21335
rect 20269 21301 20303 21335
rect 21557 21301 21591 21335
rect 22017 21301 22051 21335
rect 23305 21301 23339 21335
rect 21465 21097 21499 21131
rect 21005 21029 21039 21063
rect 10701 20961 10735 20995
rect 16957 20961 16991 20995
rect 19625 20961 19659 20995
rect 22201 20961 22235 20995
rect 24685 20961 24719 20995
rect 9965 20893 9999 20927
rect 19809 20893 19843 20927
rect 20453 20893 20487 20927
rect 20821 20893 20855 20927
rect 22661 20893 22695 20927
rect 23857 20893 23891 20927
rect 10977 20825 11011 20859
rect 16681 20825 16715 20859
rect 19717 20825 19751 20859
rect 21281 20825 21315 20859
rect 9137 20757 9171 20791
rect 12449 20757 12483 20791
rect 12725 20757 12759 20791
rect 14657 20757 14691 20791
rect 15209 20757 15243 20791
rect 17233 20757 17267 20791
rect 18705 20757 18739 20791
rect 20177 20757 20211 20791
rect 24869 20757 24903 20791
rect 24961 20757 24995 20791
rect 25329 20757 25363 20791
rect 10057 20553 10091 20587
rect 10425 20553 10459 20587
rect 10793 20553 10827 20587
rect 15301 20553 15335 20587
rect 23305 20553 23339 20587
rect 25329 20553 25363 20587
rect 20821 20485 20855 20519
rect 21465 20485 21499 20519
rect 7757 20417 7791 20451
rect 12725 20417 12759 20451
rect 15393 20417 15427 20451
rect 18613 20417 18647 20451
rect 19257 20417 19291 20451
rect 19901 20417 19935 20451
rect 22017 20417 22051 20451
rect 22753 20417 22787 20451
rect 8033 20349 8067 20383
rect 9781 20349 9815 20383
rect 10885 20349 10919 20383
rect 10977 20349 11011 20383
rect 13001 20349 13035 20383
rect 15117 20349 15151 20383
rect 18337 20349 18371 20383
rect 20545 20349 20579 20383
rect 20729 20349 20763 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 22201 20281 22235 20315
rect 14473 20213 14507 20247
rect 15761 20213 15795 20247
rect 16865 20213 16899 20247
rect 19073 20213 19107 20247
rect 19717 20213 19751 20247
rect 21189 20213 21223 20247
rect 22937 20213 22971 20247
rect 10885 20009 10919 20043
rect 12081 20009 12115 20043
rect 16037 20009 16071 20043
rect 16681 20009 16715 20043
rect 18245 20009 18279 20043
rect 23857 20009 23891 20043
rect 16957 19941 16991 19975
rect 9413 19873 9447 19907
rect 11529 19873 11563 19907
rect 14289 19873 14323 19907
rect 17693 19873 17727 19907
rect 19901 19873 19935 19907
rect 22109 19873 22143 19907
rect 9137 19805 9171 19839
rect 16497 19805 16531 19839
rect 17785 19805 17819 19839
rect 18889 19805 18923 19839
rect 14565 19737 14599 19771
rect 17877 19737 17911 19771
rect 20177 19737 20211 19771
rect 22385 19737 22419 19771
rect 24133 19737 24167 19771
rect 24409 19737 24443 19771
rect 24593 19737 24627 19771
rect 8401 19669 8435 19703
rect 11621 19669 11655 19703
rect 11713 19669 11747 19703
rect 18705 19669 18739 19703
rect 21649 19669 21683 19703
rect 24869 19669 24903 19703
rect 8769 19465 8803 19499
rect 10977 19465 11011 19499
rect 11713 19465 11747 19499
rect 12541 19465 12575 19499
rect 15209 19465 15243 19499
rect 17141 19465 17175 19499
rect 17601 19465 17635 19499
rect 20453 19465 20487 19499
rect 20545 19465 20579 19499
rect 22201 19465 22235 19499
rect 22661 19465 22695 19499
rect 25145 19465 25179 19499
rect 14013 19397 14047 19431
rect 23673 19397 23707 19431
rect 9137 19329 9171 19363
rect 9229 19329 9263 19363
rect 14289 19329 14323 19363
rect 15025 19329 15059 19363
rect 16129 19329 16163 19363
rect 17233 19329 17267 19363
rect 18981 19329 19015 19363
rect 21465 19329 21499 19363
rect 22569 19329 22603 19363
rect 23397 19329 23431 19363
rect 6561 19261 6595 19295
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 16957 19261 16991 19295
rect 20729 19261 20763 19295
rect 22845 19261 22879 19295
rect 11253 19193 11287 19227
rect 15945 19193 15979 19227
rect 8309 19125 8343 19159
rect 14565 19125 14599 19159
rect 19165 19125 19199 19159
rect 20085 19125 20119 19159
rect 21833 19125 21867 19159
rect 8401 18921 8435 18955
rect 10793 18921 10827 18955
rect 12265 18921 12299 18955
rect 17877 18921 17911 18955
rect 25237 18921 25271 18955
rect 12725 18853 12759 18887
rect 6929 18785 6963 18819
rect 10241 18785 10275 18819
rect 11621 18785 11655 18819
rect 11805 18785 11839 18819
rect 13277 18785 13311 18819
rect 16957 18785 16991 18819
rect 23857 18785 23891 18819
rect 6653 18717 6687 18751
rect 17233 18717 17267 18751
rect 21465 18717 21499 18751
rect 22017 18717 22051 18751
rect 22753 18717 22787 18751
rect 24777 18717 24811 18751
rect 8677 18649 8711 18683
rect 10425 18649 10459 18683
rect 11069 18649 11103 18683
rect 11897 18649 11931 18683
rect 18061 18649 18095 18683
rect 9689 18581 9723 18615
rect 10333 18581 10367 18615
rect 13093 18581 13127 18615
rect 13185 18581 13219 18615
rect 13829 18581 13863 18615
rect 14289 18581 14323 18615
rect 17141 18581 17175 18615
rect 17601 18581 17635 18615
rect 21281 18581 21315 18615
rect 22201 18581 22235 18615
rect 24685 18581 24719 18615
rect 13829 18377 13863 18411
rect 14289 18377 14323 18411
rect 14933 18377 14967 18411
rect 10241 18309 10275 18343
rect 13277 18309 13311 18343
rect 23305 18309 23339 18343
rect 9505 18241 9539 18275
rect 10333 18241 10367 18275
rect 11069 18241 11103 18275
rect 12449 18241 12483 18275
rect 14197 18241 14231 18275
rect 16865 18241 16899 18275
rect 21281 18241 21315 18275
rect 22201 18241 22235 18275
rect 23949 18241 23983 18275
rect 7757 18173 7791 18207
rect 9229 18173 9263 18207
rect 10057 18173 10091 18207
rect 11253 18173 11287 18207
rect 14381 18173 14415 18207
rect 17141 18173 17175 18207
rect 24593 18173 24627 18207
rect 10701 18105 10735 18139
rect 18613 18037 18647 18071
rect 18981 18037 19015 18071
rect 21097 18037 21131 18071
rect 8585 17833 8619 17867
rect 13001 17833 13035 17867
rect 18429 17833 18463 17867
rect 14197 17765 14231 17799
rect 21465 17765 21499 17799
rect 7941 17697 7975 17731
rect 9781 17697 9815 17731
rect 10057 17697 10091 17731
rect 12449 17697 12483 17731
rect 16957 17697 16991 17731
rect 17969 17697 18003 17731
rect 19533 17697 19567 17731
rect 23305 17697 23339 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 8125 17629 8159 17663
rect 11805 17629 11839 17663
rect 12633 17629 12667 17663
rect 16681 17629 16715 17663
rect 17785 17629 17819 17663
rect 18797 17629 18831 17663
rect 19717 17629 19751 17663
rect 20637 17629 20671 17663
rect 21281 17629 21315 17663
rect 21925 17629 21959 17663
rect 22109 17629 22143 17663
rect 23857 17629 23891 17663
rect 8217 17561 8251 17595
rect 12541 17561 12575 17595
rect 7389 17493 7423 17527
rect 9321 17493 9355 17527
rect 13461 17493 13495 17527
rect 15669 17493 15703 17527
rect 17417 17493 17451 17527
rect 17877 17493 17911 17527
rect 18613 17493 18647 17527
rect 19809 17493 19843 17527
rect 20177 17493 20211 17527
rect 20821 17493 20855 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 8033 17289 8067 17323
rect 9413 17289 9447 17323
rect 9781 17289 9815 17323
rect 11621 17289 11655 17323
rect 11989 17289 12023 17323
rect 13185 17289 13219 17323
rect 13553 17289 13587 17323
rect 20361 17289 20395 17323
rect 22017 17289 22051 17323
rect 22753 17289 22787 17323
rect 10333 17221 10367 17255
rect 11161 17221 11195 17255
rect 17049 17221 17083 17255
rect 18061 17221 18095 17255
rect 18889 17221 18923 17255
rect 20637 17221 20671 17255
rect 23765 17221 23799 17255
rect 7389 17153 7423 17187
rect 7941 17153 7975 17187
rect 8769 17153 8803 17187
rect 9321 17153 9355 17187
rect 16313 17153 16347 17187
rect 21465 17153 21499 17187
rect 22661 17153 22695 17187
rect 23489 17153 23523 17187
rect 7849 17085 7883 17119
rect 9229 17085 9263 17119
rect 12909 17085 12943 17119
rect 13093 17085 13127 17119
rect 14565 17085 14599 17119
rect 16037 17085 16071 17119
rect 17877 17085 17911 17119
rect 18613 17085 18647 17119
rect 22937 17085 22971 17119
rect 25237 17085 25271 17119
rect 12081 17017 12115 17051
rect 12541 17017 12575 17051
rect 8401 16949 8435 16983
rect 16957 16949 16991 16983
rect 17509 16949 17543 16983
rect 22293 16949 22327 16983
rect 8493 16745 8527 16779
rect 13921 16745 13955 16779
rect 22293 16745 22327 16779
rect 24593 16745 24627 16779
rect 11253 16677 11287 16711
rect 10425 16609 10459 16643
rect 10517 16609 10551 16643
rect 13277 16609 13311 16643
rect 13553 16609 13587 16643
rect 14657 16609 14691 16643
rect 15853 16609 15887 16643
rect 17969 16609 18003 16643
rect 20269 16609 20303 16643
rect 20545 16609 20579 16643
rect 22017 16609 22051 16643
rect 16129 16541 16163 16575
rect 18705 16541 18739 16575
rect 19809 16541 19843 16575
rect 22661 16541 22695 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 17233 16473 17267 16507
rect 19257 16473 19291 16507
rect 9873 16405 9907 16439
rect 10609 16405 10643 16439
rect 10977 16405 11011 16439
rect 11805 16405 11839 16439
rect 14197 16405 14231 16439
rect 14841 16405 14875 16439
rect 14933 16405 14967 16439
rect 15301 16405 15335 16439
rect 16037 16405 16071 16439
rect 16497 16405 16531 16439
rect 16865 16405 16899 16439
rect 18889 16405 18923 16439
rect 19625 16405 19659 16439
rect 11897 16201 11931 16235
rect 12173 16201 12207 16235
rect 13369 16201 13403 16235
rect 13737 16201 13771 16235
rect 14565 16201 14599 16235
rect 15761 16201 15795 16235
rect 16773 16201 16807 16235
rect 17325 16133 17359 16167
rect 19257 16133 19291 16167
rect 20085 16133 20119 16167
rect 21005 16133 21039 16167
rect 22293 16133 22327 16167
rect 6561 16065 6595 16099
rect 12541 16065 12575 16099
rect 14933 16065 14967 16099
rect 18061 16065 18095 16099
rect 18705 16065 18739 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 24777 16065 24811 16099
rect 6837 15997 6871 16031
rect 12633 15997 12667 16031
rect 12725 15997 12759 16031
rect 13829 15997 13863 16031
rect 13921 15997 13955 16031
rect 15025 15997 15059 16031
rect 15117 15997 15151 16031
rect 20913 15997 20947 16031
rect 24041 15997 24075 16031
rect 24501 15997 24535 16031
rect 17877 15929 17911 15963
rect 8309 15861 8343 15895
rect 8585 15861 8619 15895
rect 16221 15861 16255 15895
rect 17233 15861 17267 15895
rect 18521 15861 18555 15895
rect 21465 15861 21499 15895
rect 23765 15861 23799 15895
rect 9137 15657 9171 15691
rect 11621 15657 11655 15691
rect 16405 15657 16439 15691
rect 15485 15589 15519 15623
rect 21833 15589 21867 15623
rect 25053 15589 25087 15623
rect 25237 15589 25271 15623
rect 9689 15521 9723 15555
rect 12173 15521 12207 15555
rect 12633 15521 12667 15555
rect 18153 15521 18187 15555
rect 19441 15521 19475 15555
rect 22293 15521 22327 15555
rect 24041 15521 24075 15555
rect 24777 15521 24811 15555
rect 9597 15453 9631 15487
rect 10241 15453 10275 15487
rect 21649 15453 21683 15487
rect 11989 15385 12023 15419
rect 17877 15385 17911 15419
rect 19717 15385 19751 15419
rect 23765 15385 23799 15419
rect 9505 15317 9539 15351
rect 12081 15317 12115 15351
rect 13277 15317 13311 15351
rect 14289 15317 14323 15351
rect 14749 15317 14783 15351
rect 15945 15317 15979 15351
rect 18521 15317 18555 15351
rect 21189 15317 21223 15351
rect 10149 15113 10183 15147
rect 11345 15113 11379 15147
rect 12173 15113 12207 15147
rect 14105 15113 14139 15147
rect 14473 15113 14507 15147
rect 15945 15113 15979 15147
rect 16313 15113 16347 15147
rect 17509 15113 17543 15147
rect 19901 15113 19935 15147
rect 20821 15113 20855 15147
rect 18797 15045 18831 15079
rect 23305 15045 23339 15079
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 14013 14977 14047 15011
rect 19993 14977 20027 15011
rect 21005 14977 21039 15011
rect 21281 14977 21315 15011
rect 22109 14977 22143 15011
rect 24133 14977 24167 15011
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 9689 14909 9723 14943
rect 10701 14909 10735 14943
rect 13369 14909 13403 14943
rect 13921 14909 13955 14943
rect 15761 14909 15795 14943
rect 15853 14909 15887 14943
rect 19809 14909 19843 14943
rect 24685 14909 24719 14943
rect 18613 14841 18647 14875
rect 20361 14841 20395 14875
rect 12541 14773 12575 14807
rect 15301 14773 15335 14807
rect 8217 14569 8251 14603
rect 13185 14569 13219 14603
rect 15393 14501 15427 14535
rect 6469 14433 6503 14467
rect 6745 14433 6779 14467
rect 11989 14433 12023 14467
rect 12541 14433 12575 14467
rect 13553 14433 13587 14467
rect 14933 14433 14967 14467
rect 16589 14433 16623 14467
rect 21649 14433 21683 14467
rect 21741 14433 21775 14467
rect 23397 14433 23431 14467
rect 9965 14365 9999 14399
rect 14749 14365 14783 14399
rect 20453 14365 20487 14399
rect 24041 14365 24075 14399
rect 25053 14365 25087 14399
rect 10241 14297 10275 14331
rect 12725 14297 12759 14331
rect 14657 14297 14691 14331
rect 16865 14297 16899 14331
rect 17693 14297 17727 14331
rect 8585 14229 8619 14263
rect 9689 14229 9723 14263
rect 12817 14229 12851 14263
rect 13829 14229 13863 14263
rect 14289 14229 14323 14263
rect 16773 14229 16807 14263
rect 17233 14229 17267 14263
rect 20269 14229 20303 14263
rect 21833 14229 21867 14263
rect 22201 14229 22235 14263
rect 24869 14229 24903 14263
rect 12633 14025 12667 14059
rect 13001 14025 13035 14059
rect 15577 14025 15611 14059
rect 18613 14025 18647 14059
rect 19073 14025 19107 14059
rect 20361 14025 20395 14059
rect 22201 14025 22235 14059
rect 25053 14025 25087 14059
rect 11161 13957 11195 13991
rect 12265 13957 12299 13991
rect 19441 13957 19475 13991
rect 19625 13957 19659 13991
rect 7757 13889 7791 13923
rect 10333 13889 10367 13923
rect 20177 13889 20211 13923
rect 21097 13889 21131 13923
rect 22017 13889 22051 13923
rect 25237 13889 25271 13923
rect 8033 13821 8067 13855
rect 9781 13821 9815 13855
rect 11713 13821 11747 13855
rect 13093 13821 13127 13855
rect 13185 13821 13219 13855
rect 13829 13821 13863 13855
rect 15945 13821 15979 13855
rect 16865 13821 16899 13855
rect 18889 13821 18923 13855
rect 22845 13821 22879 13855
rect 24593 13821 24627 13855
rect 20913 13753 20947 13787
rect 14092 13685 14126 13719
rect 17128 13685 17162 13719
rect 23102 13685 23136 13719
rect 6561 13481 6595 13515
rect 9229 13481 9263 13515
rect 13921 13481 13955 13515
rect 17417 13481 17451 13515
rect 24593 13481 24627 13515
rect 21097 13413 21131 13447
rect 9781 13345 9815 13379
rect 12173 13345 12207 13379
rect 13461 13345 13495 13379
rect 15761 13345 15795 13379
rect 16313 13345 16347 13379
rect 23397 13345 23431 13379
rect 8309 13277 8343 13311
rect 12633 13277 12667 13311
rect 15669 13277 15703 13311
rect 17969 13277 18003 13311
rect 18705 13277 18739 13311
rect 19441 13277 19475 13311
rect 20821 13277 20855 13311
rect 21925 13277 21959 13311
rect 22201 13277 22235 13311
rect 24041 13277 24075 13311
rect 24777 13277 24811 13311
rect 8033 13209 8067 13243
rect 9597 13209 9631 13243
rect 11897 13209 11931 13243
rect 14657 13209 14691 13243
rect 15577 13209 15611 13243
rect 17785 13209 17819 13243
rect 18521 13209 18555 13243
rect 20269 13209 20303 13243
rect 25053 13209 25087 13243
rect 8677 13141 8711 13175
rect 9689 13141 9723 13175
rect 10425 13141 10459 13175
rect 14933 13141 14967 13175
rect 15209 13141 15243 13175
rect 20729 13141 20763 13175
rect 7389 12937 7423 12971
rect 9781 12937 9815 12971
rect 10793 12937 10827 12971
rect 11989 12937 12023 12971
rect 13369 12937 13403 12971
rect 14565 12937 14599 12971
rect 15025 12937 15059 12971
rect 15485 12937 15519 12971
rect 17141 12937 17175 12971
rect 17601 12937 17635 12971
rect 18245 12937 18279 12971
rect 19073 12937 19107 12971
rect 19533 12937 19567 12971
rect 22201 12937 22235 12971
rect 22753 12937 22787 12971
rect 25145 12937 25179 12971
rect 9321 12869 9355 12903
rect 10885 12869 10919 12903
rect 12081 12869 12115 12903
rect 13001 12869 13035 12903
rect 23397 12869 23431 12903
rect 7021 12801 7055 12835
rect 8125 12801 8159 12835
rect 8217 12801 8251 12835
rect 9413 12801 9447 12835
rect 11621 12801 11655 12835
rect 14197 12801 14231 12835
rect 15393 12801 15427 12835
rect 17233 12801 17267 12835
rect 18061 12801 18095 12835
rect 19165 12801 19199 12835
rect 20177 12801 20211 12835
rect 21097 12801 21131 12835
rect 22017 12801 22051 12835
rect 23121 12801 23155 12835
rect 6837 12733 6871 12767
rect 6929 12733 6963 12767
rect 8033 12733 8067 12767
rect 9137 12733 9171 12767
rect 10977 12733 11011 12767
rect 12725 12733 12759 12767
rect 12909 12733 12943 12767
rect 14013 12733 14047 12767
rect 14105 12733 14139 12767
rect 15577 12733 15611 12767
rect 17049 12733 17083 12767
rect 18981 12733 19015 12767
rect 20913 12733 20947 12767
rect 21005 12733 21039 12767
rect 22477 12733 22511 12767
rect 10425 12665 10459 12699
rect 11713 12665 11747 12699
rect 16129 12665 16163 12699
rect 8585 12597 8619 12631
rect 12265 12597 12299 12631
rect 19993 12597 20027 12631
rect 21465 12597 21499 12631
rect 24869 12597 24903 12631
rect 10241 12393 10275 12427
rect 11437 12393 11471 12427
rect 12633 12393 12667 12427
rect 14289 12393 14323 12427
rect 15301 12393 15335 12427
rect 24593 12393 24627 12427
rect 13645 12325 13679 12359
rect 15485 12325 15519 12359
rect 19993 12325 20027 12359
rect 7389 12257 7423 12291
rect 8217 12257 8251 12291
rect 10701 12257 10735 12291
rect 10793 12257 10827 12291
rect 12081 12257 12115 12291
rect 13093 12257 13127 12291
rect 13277 12257 13311 12291
rect 13921 12257 13955 12291
rect 14749 12257 14783 12291
rect 14841 12257 14875 12291
rect 18889 12257 18923 12291
rect 21925 12257 21959 12291
rect 23397 12257 23431 12291
rect 11805 12189 11839 12223
rect 16405 12189 16439 12223
rect 18245 12189 18279 12223
rect 19533 12189 19567 12223
rect 22201 12189 22235 12223
rect 24041 12189 24075 12223
rect 24777 12189 24811 12223
rect 10609 12121 10643 12155
rect 17417 12121 17451 12155
rect 19717 12121 19751 12155
rect 8953 12053 8987 12087
rect 11897 12053 11931 12087
rect 13001 12053 13035 12087
rect 14657 12053 14691 12087
rect 15669 12053 15703 12087
rect 16865 12053 16899 12087
rect 20453 12053 20487 12087
rect 7297 11849 7331 11883
rect 9873 11849 9907 11883
rect 10241 11849 10275 11883
rect 12173 11849 12207 11883
rect 12633 11849 12667 11883
rect 14289 11849 14323 11883
rect 17141 11849 17175 11883
rect 18337 11849 18371 11883
rect 18429 11849 18463 11883
rect 18797 11849 18831 11883
rect 21189 11849 21223 11883
rect 21465 11849 21499 11883
rect 8769 11781 8803 11815
rect 10333 11781 10367 11815
rect 20085 11781 20119 11815
rect 21557 11781 21591 11815
rect 11621 11713 11655 11747
rect 12265 11713 12299 11747
rect 13461 11713 13495 11747
rect 14657 11713 14691 11747
rect 15301 11713 15335 11747
rect 15577 11713 15611 11747
rect 17233 11713 17267 11747
rect 19349 11713 19383 11747
rect 23489 11713 23523 11747
rect 25145 11713 25179 11747
rect 9045 11645 9079 11679
rect 10425 11645 10459 11679
rect 11989 11645 12023 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 14749 11645 14783 11679
rect 14841 11645 14875 11679
rect 16957 11645 16991 11679
rect 18245 11645 18279 11679
rect 20729 11645 20763 11679
rect 23029 11645 23063 11679
rect 24777 11645 24811 11679
rect 9505 11577 9539 11611
rect 13093 11577 13127 11611
rect 17601 11577 17635 11611
rect 9413 11509 9447 11543
rect 11345 11509 11379 11543
rect 19441 11509 19475 11543
rect 20177 11509 20211 11543
rect 17233 11305 17267 11339
rect 17877 11305 17911 11339
rect 20361 11305 20395 11339
rect 22109 11305 22143 11339
rect 25053 11305 25087 11339
rect 10885 11237 10919 11271
rect 12173 11237 12207 11271
rect 13737 11237 13771 11271
rect 16681 11237 16715 11271
rect 18889 11237 18923 11271
rect 9413 11169 9447 11203
rect 11529 11169 11563 11203
rect 11713 11169 11747 11203
rect 13185 11169 13219 11203
rect 13829 11169 13863 11203
rect 14933 11169 14967 11203
rect 18337 11169 18371 11203
rect 19809 11169 19843 11203
rect 23305 11169 23339 11203
rect 9137 11101 9171 11135
rect 13093 11101 13127 11135
rect 18429 11101 18463 11135
rect 19257 11101 19291 11135
rect 19993 11101 20027 11135
rect 21005 11101 21039 11135
rect 21557 11101 21591 11135
rect 24041 11101 24075 11135
rect 25237 11101 25271 11135
rect 14289 11033 14323 11067
rect 15209 11033 15243 11067
rect 16957 11033 16991 11067
rect 17601 11033 17635 11067
rect 18521 11033 18555 11067
rect 20821 11033 20855 11067
rect 11805 10965 11839 10999
rect 12633 10965 12667 10999
rect 13001 10965 13035 10999
rect 19901 10965 19935 10999
rect 21741 10965 21775 10999
rect 9965 10761 9999 10795
rect 12633 10761 12667 10795
rect 12725 10761 12759 10795
rect 13829 10761 13863 10795
rect 15577 10761 15611 10795
rect 15945 10761 15979 10795
rect 17049 10761 17083 10795
rect 20269 10761 20303 10795
rect 8493 10693 8527 10727
rect 23397 10693 23431 10727
rect 25145 10693 25179 10727
rect 14197 10625 14231 10659
rect 16865 10625 16899 10659
rect 17693 10625 17727 10659
rect 18245 10625 18279 10659
rect 19073 10625 19107 10659
rect 19901 10625 19935 10659
rect 21097 10625 21131 10659
rect 22201 10625 22235 10659
rect 8217 10557 8251 10591
rect 11253 10557 11287 10591
rect 11897 10557 11931 10591
rect 12449 10557 12483 10591
rect 14289 10557 14323 10591
rect 14381 10557 14415 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 19625 10557 19659 10591
rect 19809 10557 19843 10591
rect 21189 10557 21223 10591
rect 21281 10557 21315 10591
rect 23121 10557 23155 10591
rect 13461 10489 13495 10523
rect 17509 10489 17543 10523
rect 18429 10489 18463 10523
rect 20729 10489 20763 10523
rect 7849 10421 7883 10455
rect 10425 10421 10459 10455
rect 10977 10421 11011 10455
rect 13093 10421 13127 10455
rect 15301 10421 15335 10455
rect 18889 10421 18923 10455
rect 22017 10421 22051 10455
rect 22477 10421 22511 10455
rect 22753 10421 22787 10455
rect 24869 10421 24903 10455
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 14565 10217 14599 10251
rect 15577 10217 15611 10251
rect 20177 10217 20211 10251
rect 24593 10217 24627 10251
rect 12817 10149 12851 10183
rect 9321 10081 9355 10115
rect 12173 10081 12207 10115
rect 13461 10081 13495 10115
rect 14289 10081 14323 10115
rect 15117 10081 15151 10115
rect 18429 10081 18463 10115
rect 18613 10081 18647 10115
rect 20821 10081 20855 10115
rect 23305 10081 23339 10115
rect 23397 10081 23431 10115
rect 13185 10013 13219 10047
rect 16865 10013 16899 10047
rect 20545 10013 20579 10047
rect 24777 10013 24811 10047
rect 9597 9945 9631 9979
rect 11989 9945 12023 9979
rect 13921 9945 13955 9979
rect 15025 9945 15059 9979
rect 18337 9945 18371 9979
rect 19073 9945 19107 9979
rect 19625 9945 19659 9979
rect 12081 9877 12115 9911
rect 13277 9877 13311 9911
rect 14933 9877 14967 9911
rect 15853 9877 15887 9911
rect 16313 9877 16347 9911
rect 16957 9877 16991 9911
rect 17969 9877 18003 9911
rect 19533 9877 19567 9911
rect 19993 9877 20027 9911
rect 22293 9877 22327 9911
rect 22845 9877 22879 9911
rect 23213 9877 23247 9911
rect 22017 9673 22051 9707
rect 25329 9673 25363 9707
rect 18797 9605 18831 9639
rect 24133 9605 24167 9639
rect 14289 9537 14323 9571
rect 15485 9537 15519 9571
rect 19073 9537 19107 9571
rect 20085 9537 20119 9571
rect 21281 9537 21315 9571
rect 25053 9537 25087 9571
rect 11713 9469 11747 9503
rect 11989 9469 12023 9503
rect 13461 9469 13495 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 15577 9469 15611 9503
rect 15761 9469 15795 9503
rect 16957 9469 16991 9503
rect 22661 9469 22695 9503
rect 24409 9469 24443 9503
rect 13921 9401 13955 9435
rect 15117 9401 15151 9435
rect 17325 9401 17359 9435
rect 19441 9401 19475 9435
rect 11345 9333 11379 9367
rect 16129 9333 16163 9367
rect 16405 9333 16439 9367
rect 16865 9333 16899 9367
rect 24869 9333 24903 9367
rect 14289 9129 14323 9163
rect 15945 9129 15979 9163
rect 19625 9129 19659 9163
rect 13001 9061 13035 9095
rect 15485 9061 15519 9095
rect 17141 9061 17175 9095
rect 10609 8993 10643 9027
rect 13553 8993 13587 9027
rect 14841 8993 14875 9027
rect 16497 8993 16531 9027
rect 17693 8993 17727 9027
rect 21373 8993 21407 9027
rect 25053 8993 25087 9027
rect 10885 8925 10919 8959
rect 12725 8925 12759 8959
rect 17601 8925 17635 8959
rect 18705 8925 18739 8959
rect 22017 8925 22051 8959
rect 22845 8925 22879 8959
rect 24593 8925 24627 8959
rect 13369 8857 13403 8891
rect 14749 8857 14783 8891
rect 16405 8857 16439 8891
rect 17509 8857 17543 8891
rect 18889 8857 18923 8891
rect 21097 8857 21131 8891
rect 23857 8857 23891 8891
rect 9137 8789 9171 8823
rect 11253 8789 11287 8823
rect 13461 8789 13495 8823
rect 14657 8789 14691 8823
rect 15393 8789 15427 8823
rect 16313 8789 16347 8823
rect 18245 8789 18279 8823
rect 21833 8789 21867 8823
rect 22385 8789 22419 8823
rect 24777 8789 24811 8823
rect 12909 8585 12943 8619
rect 13921 8517 13955 8551
rect 14473 8517 14507 8551
rect 25145 8517 25179 8551
rect 15393 8449 15427 8483
rect 17233 8449 17267 8483
rect 17877 8449 17911 8483
rect 18429 8449 18463 8483
rect 21465 8449 21499 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 11713 8381 11747 8415
rect 13369 8381 13403 8415
rect 15669 8381 15703 8415
rect 16129 8381 16163 8415
rect 17049 8381 17083 8415
rect 17141 8381 17175 8415
rect 19073 8381 19107 8415
rect 20453 8381 20487 8415
rect 22569 8381 22603 8415
rect 14105 8313 14139 8347
rect 17601 8313 17635 8347
rect 15853 8041 15887 8075
rect 11805 7973 11839 8007
rect 15025 7973 15059 8007
rect 23857 7973 23891 8007
rect 24593 7973 24627 8007
rect 11253 7905 11287 7939
rect 13185 7905 13219 7939
rect 14381 7905 14415 7939
rect 16405 7905 16439 7939
rect 18429 7905 18463 7939
rect 21189 7905 21223 7939
rect 22385 7905 22419 7939
rect 11437 7837 11471 7871
rect 13369 7837 13403 7871
rect 14657 7837 14691 7871
rect 18889 7837 18923 7871
rect 21649 7837 21683 7871
rect 22109 7837 22143 7871
rect 13277 7769 13311 7803
rect 16313 7769 16347 7803
rect 24777 7769 24811 7803
rect 11345 7701 11379 7735
rect 12541 7701 12575 7735
rect 13737 7701 13771 7735
rect 14565 7701 14599 7735
rect 15393 7701 15427 7735
rect 16221 7701 16255 7735
rect 19441 7701 19475 7735
rect 19901 7701 19935 7735
rect 24225 7701 24259 7735
rect 11897 7497 11931 7531
rect 12633 7497 12667 7531
rect 13001 7497 13035 7531
rect 17785 7497 17819 7531
rect 18521 7497 18555 7531
rect 21189 7497 21223 7531
rect 15209 7429 15243 7463
rect 16773 7429 16807 7463
rect 25145 7429 25179 7463
rect 9045 7361 9079 7395
rect 16129 7361 16163 7395
rect 17693 7361 17727 7395
rect 20269 7361 20303 7395
rect 21097 7361 21131 7395
rect 23305 7361 23339 7395
rect 24041 7361 24075 7395
rect 9321 7293 9355 7327
rect 12357 7293 12391 7327
rect 12541 7293 12575 7327
rect 15485 7293 15519 7327
rect 16865 7293 16899 7327
rect 17969 7293 18003 7327
rect 19993 7293 20027 7327
rect 21281 7293 21315 7327
rect 23029 7293 23063 7327
rect 11161 7225 11195 7259
rect 16313 7225 16347 7259
rect 10793 7157 10827 7191
rect 11345 7157 11379 7191
rect 13737 7157 13771 7191
rect 17325 7157 17359 7191
rect 20729 7157 20763 7191
rect 20453 6885 20487 6919
rect 12541 6817 12575 6851
rect 12909 6817 12943 6851
rect 17141 6817 17175 6851
rect 18889 6817 18923 6851
rect 19625 6817 19659 6851
rect 21741 6817 21775 6851
rect 25053 6817 25087 6851
rect 25145 6817 25179 6851
rect 10793 6749 10827 6783
rect 13553 6749 13587 6783
rect 14565 6749 14599 6783
rect 16681 6749 16715 6783
rect 22017 6749 22051 6783
rect 22661 6749 22695 6783
rect 11069 6681 11103 6715
rect 14749 6681 14783 6715
rect 15761 6681 15795 6715
rect 17417 6681 17451 6715
rect 19809 6681 19843 6715
rect 23857 6681 23891 6715
rect 24961 6681 24995 6715
rect 13737 6613 13771 6647
rect 14289 6613 14323 6647
rect 19717 6613 19751 6647
rect 20177 6613 20211 6647
rect 24593 6613 24627 6647
rect 11989 6409 12023 6443
rect 12817 6409 12851 6443
rect 14105 6409 14139 6443
rect 17325 6409 17359 6443
rect 17969 6409 18003 6443
rect 22017 6409 22051 6443
rect 24593 6409 24627 6443
rect 25053 6409 25087 6443
rect 10701 6341 10735 6375
rect 20545 6341 20579 6375
rect 10793 6273 10827 6307
rect 12081 6273 12115 6307
rect 13737 6273 13771 6307
rect 16313 6273 16347 6307
rect 17233 6273 17267 6307
rect 18245 6273 18279 6307
rect 19441 6273 19475 6307
rect 21465 6273 21499 6307
rect 23765 6273 23799 6307
rect 24777 6273 24811 6307
rect 10517 6205 10551 6239
rect 11805 6205 11839 6239
rect 13553 6205 13587 6239
rect 13645 6205 13679 6239
rect 14381 6205 14415 6239
rect 15853 6205 15887 6239
rect 17417 6205 17451 6239
rect 23489 6205 23523 6239
rect 24041 6205 24075 6239
rect 11161 6137 11195 6171
rect 16865 6137 16899 6171
rect 12449 6069 12483 6103
rect 13001 6069 13035 6103
rect 24225 6069 24259 6103
rect 25237 6069 25271 6103
rect 11805 5865 11839 5899
rect 13737 5865 13771 5899
rect 16208 5865 16242 5899
rect 17693 5865 17727 5899
rect 23857 5865 23891 5899
rect 13093 5797 13127 5831
rect 15485 5797 15519 5831
rect 24593 5797 24627 5831
rect 10333 5729 10367 5763
rect 14933 5729 14967 5763
rect 18613 5729 18647 5763
rect 18705 5729 18739 5763
rect 10057 5661 10091 5695
rect 12265 5661 12299 5695
rect 12909 5661 12943 5695
rect 13553 5661 13587 5695
rect 15117 5661 15151 5695
rect 15945 5661 15979 5695
rect 18521 5661 18555 5695
rect 20821 5661 20855 5695
rect 22477 5661 22511 5695
rect 23213 5661 23247 5695
rect 24041 5661 24075 5695
rect 24777 5661 24811 5695
rect 14473 5593 14507 5627
rect 19625 5593 19659 5627
rect 21465 5593 21499 5627
rect 23397 5593 23431 5627
rect 12449 5525 12483 5559
rect 14289 5525 14323 5559
rect 15025 5525 15059 5559
rect 18153 5525 18187 5559
rect 10057 5253 10091 5287
rect 13461 5253 13495 5287
rect 21005 5253 21039 5287
rect 21557 5253 21591 5287
rect 10333 5185 10367 5219
rect 11161 5185 11195 5219
rect 12265 5185 12299 5219
rect 12909 5185 12943 5219
rect 13185 5185 13219 5219
rect 15485 5185 15519 5219
rect 18337 5185 18371 5219
rect 20545 5185 20579 5219
rect 21189 5185 21223 5219
rect 22109 5185 22143 5219
rect 23857 5185 23891 5219
rect 12541 5117 12575 5151
rect 15761 5117 15795 5151
rect 17877 5117 17911 5151
rect 18797 5117 18831 5151
rect 20269 5117 20303 5151
rect 22477 5117 22511 5151
rect 24317 5117 24351 5151
rect 10517 5049 10551 5083
rect 10977 4981 11011 5015
rect 14933 4981 14967 5015
rect 14197 4777 14231 4811
rect 16865 4777 16899 4811
rect 24133 4777 24167 4811
rect 5089 4641 5123 4675
rect 10333 4641 10367 4675
rect 10609 4641 10643 4675
rect 13277 4641 13311 4675
rect 15117 4641 15151 4675
rect 21281 4641 21315 4675
rect 24593 4641 24627 4675
rect 1593 4573 1627 4607
rect 3985 4573 4019 4607
rect 7113 4573 7147 4607
rect 11069 4573 11103 4607
rect 11345 4573 11379 4607
rect 13737 4573 13771 4607
rect 18797 4573 18831 4607
rect 21741 4573 21775 4607
rect 24777 4573 24811 4607
rect 25145 4573 25179 4607
rect 4629 4505 4663 4539
rect 5365 4505 5399 4539
rect 7389 4505 7423 4539
rect 15393 4505 15427 4539
rect 17601 4505 17635 4539
rect 21005 4505 21039 4539
rect 22661 4505 22695 4539
rect 23765 4505 23799 4539
rect 1777 4437 1811 4471
rect 9229 4437 9263 4471
rect 9505 4437 9539 4471
rect 14657 4437 14691 4471
rect 19533 4437 19567 4471
rect 23673 4437 23707 4471
rect 25329 4437 25363 4471
rect 2881 4233 2915 4267
rect 11161 4233 11195 4267
rect 15669 4233 15703 4267
rect 14197 4165 14231 4199
rect 21833 4165 21867 4199
rect 22109 4165 22143 4199
rect 22477 4165 22511 4199
rect 1593 4097 1627 4131
rect 2697 4081 2731 4115
rect 4169 4097 4203 4131
rect 4813 4097 4847 4131
rect 9045 4097 9079 4131
rect 10241 4097 10275 4131
rect 13461 4097 13495 4131
rect 13921 4097 13955 4131
rect 16313 4097 16347 4131
rect 18245 4097 18279 4131
rect 18705 4097 18739 4131
rect 20913 4097 20947 4131
rect 21005 4097 21039 4131
rect 21649 4097 21683 4131
rect 24225 4097 24259 4131
rect 24685 4097 24719 4131
rect 10517 4029 10551 4063
rect 11621 4029 11655 4063
rect 13001 4029 13035 4063
rect 17049 4029 17083 4063
rect 19165 4029 19199 4063
rect 21097 4029 21131 4063
rect 3249 3961 3283 3995
rect 4353 3961 4387 3995
rect 5365 3961 5399 3995
rect 7113 3961 7147 3995
rect 16129 3961 16163 3995
rect 2237 3893 2271 3927
rect 3433 3893 3467 3927
rect 3893 3893 3927 3927
rect 4997 3893 5031 3927
rect 6101 3893 6135 3927
rect 7021 3893 7055 3927
rect 7481 3893 7515 3927
rect 7757 3893 7791 3927
rect 8033 3893 8067 3927
rect 9229 3893 9263 3927
rect 11805 3893 11839 3927
rect 20545 3893 20579 3927
rect 25329 3893 25363 3927
rect 1961 3689 1995 3723
rect 4445 3689 4479 3723
rect 8585 3689 8619 3723
rect 9873 3689 9907 3723
rect 18659 3689 18693 3723
rect 24041 3689 24075 3723
rect 3249 3621 3283 3655
rect 10609 3621 10643 3655
rect 3985 3553 4019 3587
rect 4905 3553 4939 3587
rect 5181 3553 5215 3587
rect 11621 3553 11655 3587
rect 19901 3553 19935 3587
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 4261 3485 4295 3519
rect 6377 3485 6411 3519
rect 7113 3485 7147 3519
rect 7757 3485 7791 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9689 3485 9723 3519
rect 10425 3485 10459 3519
rect 11897 3485 11931 3519
rect 13737 3485 13771 3519
rect 15669 3485 15703 3519
rect 17509 3485 17543 3519
rect 18889 3485 18923 3519
rect 19533 3485 19567 3519
rect 21281 3485 21315 3519
rect 22201 3485 22235 3519
rect 23397 3485 23431 3519
rect 25237 3485 25271 3519
rect 9413 3417 9447 3451
rect 12817 3417 12851 3451
rect 14473 3417 14507 3451
rect 16313 3417 16347 3451
rect 1501 3349 1535 3383
rect 6101 3349 6135 3383
rect 6561 3349 6595 3383
rect 7297 3349 7331 3383
rect 7941 3349 7975 3383
rect 22937 3349 22971 3383
rect 24593 3349 24627 3383
rect 4537 3145 4571 3179
rect 6745 3145 6779 3179
rect 9873 3145 9907 3179
rect 11161 3145 11195 3179
rect 21281 3145 21315 3179
rect 22201 3145 22235 3179
rect 23581 3145 23615 3179
rect 25053 3145 25087 3179
rect 9413 3077 9447 3111
rect 18889 3077 18923 3111
rect 20637 3077 20671 3111
rect 20821 3077 20855 3111
rect 22753 3077 22787 3111
rect 22937 3077 22971 3111
rect 24225 3077 24259 3111
rect 24593 3077 24627 3111
rect 25237 3077 25271 3111
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 3433 3009 3467 3043
rect 3709 3009 3743 3043
rect 6009 3009 6043 3043
rect 6561 3009 6595 3043
rect 7205 3009 7239 3043
rect 7849 3009 7883 3043
rect 8125 3009 8159 3043
rect 9045 3009 9079 3043
rect 9689 3009 9723 3043
rect 10333 3009 10367 3043
rect 10977 3009 11011 3043
rect 11989 3009 12023 3043
rect 14381 3009 14415 3043
rect 14841 3009 14875 3043
rect 18061 3009 18095 3043
rect 19901 3009 19935 3043
rect 22109 3009 22143 3043
rect 23673 3009 23707 3043
rect 25421 3009 25455 3043
rect 2421 2941 2455 2975
rect 5733 2941 5767 2975
rect 9229 2941 9263 2975
rect 11713 2941 11747 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17049 2941 17083 2975
rect 1685 2873 1719 2907
rect 10517 2873 10551 2907
rect 4905 2805 4939 2839
rect 7389 2805 7423 2839
rect 24133 2805 24167 2839
rect 4629 2601 4663 2635
rect 6837 2601 6871 2635
rect 9321 2601 9355 2635
rect 14197 2601 14231 2635
rect 16221 2601 16255 2635
rect 16405 2601 16439 2635
rect 18705 2601 18739 2635
rect 23857 2601 23891 2635
rect 7941 2533 7975 2567
rect 5457 2465 5491 2499
rect 10701 2465 10735 2499
rect 14933 2465 14967 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 21281 2465 21315 2499
rect 1685 2397 1719 2431
rect 2329 2397 2363 2431
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 5181 2397 5215 2431
rect 6469 2397 6503 2431
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 12449 2397 12483 2431
rect 14473 2397 14507 2431
rect 16865 2397 16899 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 22201 2397 22235 2431
rect 23397 2397 23431 2431
rect 24041 2397 24075 2431
rect 25237 2397 25271 2431
rect 6653 2329 6687 2363
rect 13277 2329 13311 2363
rect 1869 2261 1903 2295
rect 7297 2261 7331 2295
rect 8585 2261 8619 2295
rect 11897 2261 11931 2295
rect 24593 2261 24627 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 13814 54272 13820 54324
rect 13872 54272 13878 54324
rect 18966 54272 18972 54324
rect 19024 54272 19030 54324
rect 2406 54204 2412 54256
rect 2464 54204 2470 54256
rect 5077 54247 5135 54253
rect 5077 54213 5089 54247
rect 5123 54244 5135 54247
rect 5166 54244 5172 54256
rect 5123 54216 5172 54244
rect 5123 54213 5135 54216
rect 5077 54207 5135 54213
rect 5166 54204 5172 54216
rect 5224 54204 5230 54256
rect 3421 54179 3479 54185
rect 3421 54145 3433 54179
rect 3467 54176 3479 54179
rect 4982 54176 4988 54188
rect 3467 54148 4988 54176
rect 3467 54145 3479 54148
rect 3421 54139 3479 54145
rect 4982 54136 4988 54148
rect 5040 54136 5046 54188
rect 5994 54136 6000 54188
rect 6052 54136 6058 54188
rect 8386 54136 8392 54188
rect 8444 54136 8450 54188
rect 9582 54136 9588 54188
rect 9640 54136 9646 54188
rect 11698 54136 11704 54188
rect 11756 54176 11762 54188
rect 12161 54179 12219 54185
rect 12161 54176 12173 54179
rect 11756 54148 12173 54176
rect 11756 54136 11762 54148
rect 12161 54145 12173 54148
rect 12207 54145 12219 54179
rect 13832 54176 13860 54272
rect 14568 54216 18276 54244
rect 14461 54179 14519 54185
rect 14461 54176 14473 54179
rect 13832 54148 14473 54176
rect 12161 54139 12219 54145
rect 14461 54145 14473 54148
rect 14507 54145 14519 54179
rect 14461 54139 14519 54145
rect 7834 54068 7840 54120
rect 7892 54068 7898 54120
rect 9306 54068 9312 54120
rect 9364 54108 9370 54120
rect 9861 54111 9919 54117
rect 9861 54108 9873 54111
rect 9364 54080 9873 54108
rect 9364 54068 9370 54080
rect 9861 54077 9873 54080
rect 9907 54077 9919 54111
rect 9861 54071 9919 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12621 54111 12679 54117
rect 12621 54108 12633 54111
rect 12400 54080 12633 54108
rect 12400 54068 12406 54080
rect 12621 54077 12633 54080
rect 12667 54077 12679 54111
rect 14568 54108 14596 54216
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15105 54179 15163 54185
rect 15105 54176 15117 54179
rect 14884 54148 15117 54176
rect 14884 54136 14890 54148
rect 15105 54145 15117 54148
rect 15151 54176 15163 54179
rect 15381 54179 15439 54185
rect 15381 54176 15393 54179
rect 15151 54148 15393 54176
rect 15151 54145 15163 54148
rect 15105 54139 15163 54145
rect 15381 54145 15393 54148
rect 15427 54145 15439 54179
rect 15381 54139 15439 54145
rect 16574 54136 16580 54188
rect 16632 54176 16638 54188
rect 17037 54179 17095 54185
rect 17037 54176 17049 54179
rect 16632 54148 17049 54176
rect 16632 54136 16638 54148
rect 17037 54145 17049 54148
rect 17083 54176 17095 54179
rect 17313 54179 17371 54185
rect 17313 54176 17325 54179
rect 17083 54148 17325 54176
rect 17083 54145 17095 54148
rect 17037 54139 17095 54145
rect 17313 54145 17325 54148
rect 17359 54145 17371 54179
rect 17313 54139 17371 54145
rect 17586 54136 17592 54188
rect 17644 54176 17650 54188
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17644 54148 17877 54176
rect 17644 54136 17650 54148
rect 17865 54145 17877 54148
rect 17911 54176 17923 54179
rect 18141 54179 18199 54185
rect 18141 54176 18153 54179
rect 17911 54148 18153 54176
rect 17911 54145 17923 54148
rect 17865 54139 17923 54145
rect 18141 54145 18153 54148
rect 18187 54145 18199 54179
rect 18141 54139 18199 54145
rect 12621 54071 12679 54077
rect 12728 54080 14596 54108
rect 18248 54108 18276 54216
rect 18984 54176 19012 54272
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 18984 54148 19441 54176
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 20993 54179 21051 54185
rect 20993 54176 21005 54179
rect 20772 54148 21005 54176
rect 20772 54136 20778 54148
rect 20993 54145 21005 54148
rect 21039 54176 21051 54179
rect 21269 54179 21327 54185
rect 21269 54176 21281 54179
rect 21039 54148 21281 54176
rect 21039 54145 21051 54148
rect 20993 54139 21051 54145
rect 21269 54145 21281 54148
rect 21315 54145 21327 54179
rect 21269 54139 21327 54145
rect 22094 54136 22100 54188
rect 22152 54176 22158 54188
rect 22281 54179 22339 54185
rect 22281 54176 22293 54179
rect 22152 54148 22293 54176
rect 22152 54136 22158 54148
rect 22281 54145 22293 54148
rect 22327 54176 22339 54179
rect 22557 54179 22615 54185
rect 22557 54176 22569 54179
rect 22327 54148 22569 54176
rect 22327 54145 22339 54148
rect 22281 54139 22339 54145
rect 22557 54145 22569 54148
rect 22603 54145 22615 54179
rect 22557 54139 22615 54145
rect 24029 54179 24087 54185
rect 24029 54145 24041 54179
rect 24075 54176 24087 54179
rect 24673 54179 24731 54185
rect 24673 54176 24685 54179
rect 24075 54148 24685 54176
rect 24075 54145 24087 54148
rect 24029 54139 24087 54145
rect 24673 54145 24685 54148
rect 24719 54145 24731 54179
rect 24673 54139 24731 54145
rect 25317 54179 25375 54185
rect 25317 54145 25329 54179
rect 25363 54176 25375 54179
rect 25866 54176 25872 54188
rect 25363 54148 25872 54176
rect 25363 54145 25375 54148
rect 25317 54139 25375 54145
rect 19705 54111 19763 54117
rect 19705 54108 19717 54111
rect 18248 54080 19717 54108
rect 8478 54000 8484 54052
rect 8536 54040 8542 54052
rect 12728 54040 12756 54080
rect 19705 54077 19717 54080
rect 19751 54077 19763 54111
rect 19705 54071 19763 54077
rect 23109 54111 23167 54117
rect 23109 54077 23121 54111
rect 23155 54108 23167 54111
rect 25332 54108 25360 54139
rect 25866 54136 25872 54148
rect 25924 54136 25930 54188
rect 23155 54080 25360 54108
rect 23155 54077 23167 54080
rect 23109 54071 23167 54077
rect 8536 54012 12756 54040
rect 8536 54000 8542 54012
rect 13906 54000 13912 54052
rect 13964 54040 13970 54052
rect 14921 54043 14979 54049
rect 14921 54040 14933 54043
rect 13964 54012 14933 54040
rect 13964 54000 13970 54012
rect 14921 54009 14933 54012
rect 14967 54009 14979 54043
rect 14921 54003 14979 54009
rect 16758 54000 16764 54052
rect 16816 54040 16822 54052
rect 20809 54043 20867 54049
rect 20809 54040 20821 54043
rect 16816 54012 20821 54040
rect 16816 54000 16822 54012
rect 20809 54009 20821 54012
rect 20855 54009 20867 54043
rect 20809 54003 20867 54009
rect 12710 53932 12716 53984
rect 12768 53972 12774 53984
rect 14277 53975 14335 53981
rect 14277 53972 14289 53975
rect 12768 53944 14289 53972
rect 12768 53932 12774 53944
rect 14277 53941 14289 53944
rect 14323 53941 14335 53975
rect 14277 53935 14335 53941
rect 16850 53932 16856 53984
rect 16908 53932 16914 53984
rect 17494 53932 17500 53984
rect 17552 53972 17558 53984
rect 17681 53975 17739 53981
rect 17681 53972 17693 53975
rect 17552 53944 17693 53972
rect 17552 53932 17558 53944
rect 17681 53941 17693 53944
rect 17727 53941 17739 53975
rect 17681 53935 17739 53941
rect 22094 53932 22100 53984
rect 22152 53932 22158 53984
rect 23385 53975 23443 53981
rect 23385 53941 23397 53975
rect 23431 53972 23443 53975
rect 24670 53972 24676 53984
rect 23431 53944 24676 53972
rect 23431 53941 23443 53944
rect 23385 53935 23443 53941
rect 24670 53932 24676 53944
rect 24728 53932 24734 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 10686 53660 10692 53712
rect 10744 53660 10750 53712
rect 24854 53700 24860 53712
rect 22572 53672 24860 53700
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 1765 53635 1823 53641
rect 1765 53632 1777 53635
rect 1084 53604 1777 53632
rect 1084 53592 1090 53604
rect 1765 53601 1777 53604
rect 1811 53601 1823 53635
rect 1765 53595 1823 53601
rect 3786 53592 3792 53644
rect 3844 53632 3850 53644
rect 4157 53635 4215 53641
rect 4157 53632 4169 53635
rect 3844 53604 4169 53632
rect 3844 53592 3850 53604
rect 4157 53601 4169 53604
rect 4203 53601 4215 53635
rect 4157 53595 4215 53601
rect 6546 53592 6552 53644
rect 6604 53632 6610 53644
rect 6917 53635 6975 53641
rect 6917 53632 6929 53635
rect 6604 53604 6929 53632
rect 6604 53592 6610 53604
rect 6917 53601 6929 53604
rect 6963 53601 6975 53635
rect 10704 53632 10732 53660
rect 11241 53635 11299 53641
rect 11241 53632 11253 53635
rect 10704 53604 11253 53632
rect 6917 53595 6975 53601
rect 11241 53601 11253 53604
rect 11287 53601 11299 53635
rect 11241 53595 11299 53601
rect 22572 53576 22600 53672
rect 24854 53660 24860 53672
rect 24912 53660 24918 53712
rect 23290 53592 23296 53644
rect 23348 53632 23354 53644
rect 23348 53604 23796 53632
rect 23348 53592 23354 53604
rect 2961 53567 3019 53573
rect 2961 53533 2973 53567
rect 3007 53533 3019 53567
rect 2961 53527 3019 53533
rect 2976 53496 3004 53527
rect 5350 53524 5356 53576
rect 5408 53524 5414 53576
rect 8021 53567 8079 53573
rect 8021 53533 8033 53567
rect 8067 53564 8079 53567
rect 9214 53564 9220 53576
rect 8067 53536 9220 53564
rect 8067 53533 8079 53536
rect 8021 53527 8079 53533
rect 9214 53524 9220 53536
rect 9272 53524 9278 53576
rect 10686 53524 10692 53576
rect 10744 53564 10750 53576
rect 10781 53567 10839 53573
rect 10781 53564 10793 53567
rect 10744 53536 10793 53564
rect 10744 53524 10750 53536
rect 10781 53533 10793 53536
rect 10827 53533 10839 53567
rect 10781 53527 10839 53533
rect 22554 53524 22560 53576
rect 22612 53524 22618 53576
rect 23201 53567 23259 53573
rect 23201 53533 23213 53567
rect 23247 53564 23259 53567
rect 23382 53564 23388 53576
rect 23247 53536 23388 53564
rect 23247 53533 23259 53536
rect 23201 53527 23259 53533
rect 23382 53524 23388 53536
rect 23440 53524 23446 53576
rect 23768 53573 23796 53604
rect 23753 53567 23811 53573
rect 23753 53533 23765 53567
rect 23799 53533 23811 53567
rect 23753 53527 23811 53533
rect 24670 53524 24676 53576
rect 24728 53524 24734 53576
rect 5534 53496 5540 53508
rect 2976 53468 5540 53496
rect 5534 53456 5540 53468
rect 5592 53456 5598 53508
rect 22738 53456 22744 53508
rect 22796 53496 22802 53508
rect 23017 53499 23075 53505
rect 23017 53496 23029 53499
rect 22796 53468 23029 53496
rect 22796 53456 22802 53468
rect 23017 53465 23029 53468
rect 23063 53465 23075 53499
rect 23017 53459 23075 53465
rect 22373 53431 22431 53437
rect 22373 53397 22385 53431
rect 22419 53428 22431 53431
rect 22646 53428 22652 53440
rect 22419 53400 22652 53428
rect 22419 53397 22431 53400
rect 22373 53391 22431 53397
rect 22646 53388 22652 53400
rect 22704 53388 22710 53440
rect 23658 53388 23664 53440
rect 23716 53428 23722 53440
rect 23937 53431 23995 53437
rect 23937 53428 23949 53431
rect 23716 53400 23949 53428
rect 23716 53388 23722 53400
rect 23937 53397 23949 53400
rect 23983 53397 23995 53431
rect 23937 53391 23995 53397
rect 24578 53388 24584 53440
rect 24636 53428 24642 53440
rect 25317 53431 25375 53437
rect 25317 53428 25329 53431
rect 24636 53400 25329 53428
rect 24636 53388 24642 53400
rect 25317 53397 25329 53400
rect 25363 53397 25375 53431
rect 25317 53391 25375 53397
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 4982 53184 4988 53236
rect 5040 53224 5046 53236
rect 5169 53227 5227 53233
rect 5169 53224 5181 53227
rect 5040 53196 5181 53224
rect 5040 53184 5046 53196
rect 5169 53193 5181 53196
rect 5215 53193 5227 53227
rect 5169 53187 5227 53193
rect 22554 53184 22560 53236
rect 22612 53224 22618 53236
rect 22649 53227 22707 53233
rect 22649 53224 22661 53227
rect 22612 53196 22661 53224
rect 22612 53184 22618 53196
rect 22649 53193 22661 53196
rect 22695 53193 22707 53227
rect 22649 53187 22707 53193
rect 23290 53184 23296 53236
rect 23348 53184 23354 53236
rect 23382 53184 23388 53236
rect 23440 53184 23446 53236
rect 24762 53184 24768 53236
rect 24820 53224 24826 53236
rect 25041 53227 25099 53233
rect 25041 53224 25053 53227
rect 24820 53196 25053 53224
rect 24820 53184 24826 53196
rect 25041 53193 25053 53196
rect 25087 53193 25099 53227
rect 25041 53187 25099 53193
rect 25314 53184 25320 53236
rect 25372 53184 25378 53236
rect 24780 53156 24808 53184
rect 24044 53128 24808 53156
rect 5353 53091 5411 53097
rect 5353 53057 5365 53091
rect 5399 53088 5411 53091
rect 7558 53088 7564 53100
rect 5399 53060 7564 53088
rect 5399 53057 5411 53060
rect 5353 53051 5411 53057
rect 7558 53048 7564 53060
rect 7616 53048 7622 53100
rect 24044 53097 24072 53128
rect 24029 53091 24087 53097
rect 24029 53057 24041 53091
rect 24075 53057 24087 53091
rect 24029 53051 24087 53057
rect 24765 53091 24823 53097
rect 24765 53057 24777 53091
rect 24811 53088 24823 53091
rect 25332 53088 25360 53184
rect 24811 53060 25360 53088
rect 24811 53057 24823 53060
rect 24765 53051 24823 53057
rect 25498 52912 25504 52964
rect 25556 52912 25562 52964
rect 23842 52844 23848 52896
rect 23900 52844 23906 52896
rect 24118 52844 24124 52896
rect 24176 52884 24182 52896
rect 24581 52887 24639 52893
rect 24581 52884 24593 52887
rect 24176 52856 24593 52884
rect 24176 52844 24182 52856
rect 24581 52853 24593 52856
rect 24627 52853 24639 52887
rect 24581 52847 24639 52853
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 5350 52640 5356 52692
rect 5408 52680 5414 52692
rect 6549 52683 6607 52689
rect 6549 52680 6561 52683
rect 5408 52652 6561 52680
rect 5408 52640 5414 52652
rect 6549 52649 6561 52652
rect 6595 52649 6607 52683
rect 6549 52643 6607 52649
rect 24486 52640 24492 52692
rect 24544 52640 24550 52692
rect 23566 52572 23572 52624
rect 23624 52612 23630 52624
rect 23845 52615 23903 52621
rect 23845 52612 23857 52615
rect 23624 52584 23857 52612
rect 23624 52572 23630 52584
rect 23845 52581 23857 52584
rect 23891 52581 23903 52615
rect 23845 52575 23903 52581
rect 17402 52504 17408 52556
rect 17460 52544 17466 52556
rect 24949 52547 25007 52553
rect 24949 52544 24961 52547
rect 17460 52516 24961 52544
rect 17460 52504 17466 52516
rect 24949 52513 24961 52516
rect 24995 52513 25007 52547
rect 24949 52507 25007 52513
rect 6733 52479 6791 52485
rect 6733 52445 6745 52479
rect 6779 52476 6791 52479
rect 9398 52476 9404 52488
rect 6779 52448 9404 52476
rect 6779 52445 6791 52448
rect 6733 52439 6791 52445
rect 9398 52436 9404 52448
rect 9456 52436 9462 52488
rect 24029 52479 24087 52485
rect 24029 52445 24041 52479
rect 24075 52476 24087 52479
rect 24486 52476 24492 52488
rect 24075 52448 24492 52476
rect 24075 52445 24087 52448
rect 24029 52439 24087 52445
rect 24486 52436 24492 52448
rect 24544 52436 24550 52488
rect 25222 52368 25228 52420
rect 25280 52368 25286 52420
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 24121 52139 24179 52145
rect 24121 52105 24133 52139
rect 24167 52136 24179 52139
rect 25222 52136 25228 52148
rect 24167 52108 25228 52136
rect 24167 52105 24179 52108
rect 24121 52099 24179 52105
rect 25222 52096 25228 52108
rect 25280 52096 25286 52148
rect 24578 51960 24584 52012
rect 24636 51960 24642 52012
rect 25317 52003 25375 52009
rect 25317 51969 25329 52003
rect 25363 52000 25375 52003
rect 25498 52000 25504 52012
rect 25363 51972 25504 52000
rect 25363 51969 25375 51972
rect 25317 51963 25375 51969
rect 25498 51960 25504 51972
rect 25556 51960 25562 52012
rect 24394 51756 24400 51808
rect 24452 51756 24458 51808
rect 25133 51799 25191 51805
rect 25133 51765 25145 51799
rect 25179 51796 25191 51799
rect 26878 51796 26884 51808
rect 25179 51768 26884 51796
rect 25179 51765 25191 51768
rect 25133 51759 25191 51765
rect 26878 51756 26884 51768
rect 26936 51756 26942 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 8297 51595 8355 51601
rect 8297 51561 8309 51595
rect 8343 51592 8355 51595
rect 8386 51592 8392 51604
rect 8343 51564 8392 51592
rect 8343 51561 8355 51564
rect 8297 51555 8355 51561
rect 8386 51552 8392 51564
rect 8444 51552 8450 51604
rect 9214 51552 9220 51604
rect 9272 51552 9278 51604
rect 5994 51484 6000 51536
rect 6052 51524 6058 51536
rect 7561 51527 7619 51533
rect 7561 51524 7573 51527
rect 6052 51496 7573 51524
rect 6052 51484 6058 51496
rect 7561 51493 7573 51496
rect 7607 51493 7619 51527
rect 7561 51487 7619 51493
rect 7834 51348 7840 51400
rect 7892 51388 7898 51400
rect 8481 51391 8539 51397
rect 8481 51388 8493 51391
rect 7892 51360 8493 51388
rect 7892 51348 7898 51360
rect 8481 51357 8493 51360
rect 8527 51357 8539 51391
rect 8481 51351 8539 51357
rect 9401 51391 9459 51397
rect 9401 51357 9413 51391
rect 9447 51388 9459 51391
rect 10410 51388 10416 51400
rect 9447 51360 10416 51388
rect 9447 51357 9459 51360
rect 9401 51351 9459 51357
rect 10410 51348 10416 51360
rect 10468 51348 10474 51400
rect 7745 51323 7803 51329
rect 7745 51289 7757 51323
rect 7791 51320 7803 51323
rect 10318 51320 10324 51332
rect 7791 51292 10324 51320
rect 7791 51289 7803 51292
rect 7745 51283 7803 51289
rect 10318 51280 10324 51292
rect 10376 51280 10382 51332
rect 24581 51323 24639 51329
rect 24581 51289 24593 51323
rect 24627 51320 24639 51323
rect 25222 51320 25228 51332
rect 24627 51292 25228 51320
rect 24627 51289 24639 51292
rect 24581 51283 24639 51289
rect 25222 51280 25228 51292
rect 25280 51280 25286 51332
rect 25133 51255 25191 51261
rect 25133 51221 25145 51255
rect 25179 51252 25191 51255
rect 26510 51252 26516 51264
rect 25179 51224 26516 51252
rect 25179 51221 25191 51224
rect 25133 51215 25191 51221
rect 26510 51212 26516 51224
rect 26568 51212 26574 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 24581 50915 24639 50921
rect 24581 50881 24593 50915
rect 24627 50912 24639 50915
rect 25222 50912 25228 50924
rect 24627 50884 25228 50912
rect 24627 50881 24639 50884
rect 24581 50875 24639 50881
rect 25222 50872 25228 50884
rect 25280 50872 25286 50924
rect 25133 50711 25191 50717
rect 25133 50677 25145 50711
rect 25179 50708 25191 50711
rect 26234 50708 26240 50720
rect 25179 50680 26240 50708
rect 25179 50677 25191 50680
rect 25133 50671 25191 50677
rect 26234 50668 26240 50680
rect 26292 50668 26298 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 5534 50464 5540 50516
rect 5592 50504 5598 50516
rect 6638 50504 6644 50516
rect 5592 50476 6644 50504
rect 5592 50464 5598 50476
rect 6638 50464 6644 50476
rect 6696 50504 6702 50516
rect 7745 50507 7803 50513
rect 7745 50504 7757 50507
rect 6696 50476 7757 50504
rect 6696 50464 6702 50476
rect 7745 50473 7757 50476
rect 7791 50473 7803 50507
rect 7745 50467 7803 50473
rect 8389 50507 8447 50513
rect 8389 50473 8401 50507
rect 8435 50504 8447 50507
rect 8478 50504 8484 50516
rect 8435 50476 8484 50504
rect 8435 50473 8447 50476
rect 8389 50467 8447 50473
rect 8478 50464 8484 50476
rect 8536 50464 8542 50516
rect 9582 50464 9588 50516
rect 9640 50464 9646 50516
rect 7558 50396 7564 50448
rect 7616 50436 7622 50448
rect 9490 50436 9496 50448
rect 7616 50408 9496 50436
rect 7616 50396 7622 50408
rect 9490 50396 9496 50408
rect 9548 50396 9554 50448
rect 8021 50303 8079 50309
rect 8021 50269 8033 50303
rect 8067 50300 8079 50303
rect 8478 50300 8484 50312
rect 8067 50272 8484 50300
rect 8067 50269 8079 50272
rect 8021 50263 8079 50269
rect 8478 50260 8484 50272
rect 8536 50260 8542 50312
rect 9493 50303 9551 50309
rect 9493 50269 9505 50303
rect 9539 50300 9551 50303
rect 9582 50300 9588 50312
rect 9539 50272 9588 50300
rect 9539 50269 9551 50272
rect 9493 50263 9551 50269
rect 9582 50260 9588 50272
rect 9640 50260 9646 50312
rect 25314 50124 25320 50176
rect 25372 50164 25378 50176
rect 25409 50167 25467 50173
rect 25409 50164 25421 50167
rect 25372 50136 25421 50164
rect 25372 50124 25378 50136
rect 25409 50133 25421 50136
rect 25455 50133 25467 50167
rect 25409 50127 25467 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 25041 49759 25099 49765
rect 25041 49725 25053 49759
rect 25087 49756 25099 49759
rect 25130 49756 25136 49768
rect 25087 49728 25136 49756
rect 25087 49725 25099 49728
rect 25041 49719 25099 49725
rect 25130 49716 25136 49728
rect 25188 49716 25194 49768
rect 25314 49716 25320 49768
rect 25372 49716 25378 49768
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 10686 49308 10692 49360
rect 10744 49308 10750 49360
rect 11698 49308 11704 49360
rect 11756 49308 11762 49360
rect 10226 49104 10232 49156
rect 10284 49144 10290 49156
rect 10505 49147 10563 49153
rect 10505 49144 10517 49147
rect 10284 49116 10517 49144
rect 10284 49104 10290 49116
rect 10505 49113 10517 49116
rect 10551 49113 10563 49147
rect 10505 49107 10563 49113
rect 10962 49104 10968 49156
rect 11020 49144 11026 49156
rect 11517 49147 11575 49153
rect 11517 49144 11529 49147
rect 11020 49116 11529 49144
rect 11020 49104 11026 49116
rect 11517 49113 11529 49116
rect 11563 49113 11575 49147
rect 11517 49107 11575 49113
rect 24765 49147 24823 49153
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 25222 49144 25228 49156
rect 24811 49116 25228 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 25222 49104 25228 49116
rect 25280 49104 25286 49156
rect 25133 49079 25191 49085
rect 25133 49045 25145 49079
rect 25179 49076 25191 49079
rect 25590 49076 25596 49088
rect 25179 49048 25596 49076
rect 25179 49045 25191 49048
rect 25133 49039 25191 49045
rect 25590 49036 25596 49048
rect 25648 49036 25654 49088
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 6638 48832 6644 48884
rect 6696 48832 6702 48884
rect 8662 48804 8668 48816
rect 7682 48776 8668 48804
rect 8662 48764 8668 48776
rect 8720 48764 8726 48816
rect 8113 48671 8171 48677
rect 8113 48637 8125 48671
rect 8159 48668 8171 48671
rect 8389 48671 8447 48677
rect 8159 48640 8340 48668
rect 8159 48637 8171 48640
rect 8113 48631 8171 48637
rect 8312 48600 8340 48640
rect 8389 48637 8401 48671
rect 8435 48668 8447 48671
rect 8435 48640 8984 48668
rect 8435 48637 8447 48640
rect 8389 48631 8447 48637
rect 8846 48600 8852 48612
rect 8312 48572 8852 48600
rect 8846 48560 8852 48572
rect 8904 48560 8910 48612
rect 8662 48492 8668 48544
rect 8720 48492 8726 48544
rect 8956 48541 8984 48640
rect 8941 48535 8999 48541
rect 8941 48501 8953 48535
rect 8987 48532 8999 48535
rect 10870 48532 10876 48544
rect 8987 48504 10876 48532
rect 8987 48501 8999 48504
rect 8941 48495 8999 48501
rect 10870 48492 10876 48504
rect 10928 48492 10934 48544
rect 25222 48492 25228 48544
rect 25280 48532 25286 48544
rect 25409 48535 25467 48541
rect 25409 48532 25421 48535
rect 25280 48504 25421 48532
rect 25280 48492 25286 48504
rect 25409 48501 25421 48504
rect 25455 48501 25467 48535
rect 25409 48495 25467 48501
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 9490 48084 9496 48136
rect 9548 48124 9554 48136
rect 10356 48127 10414 48133
rect 10356 48124 10368 48127
rect 9548 48096 10368 48124
rect 9548 48084 9554 48096
rect 10356 48093 10368 48096
rect 10402 48093 10414 48127
rect 10356 48087 10414 48093
rect 24029 48127 24087 48133
rect 24029 48093 24041 48127
rect 24075 48124 24087 48127
rect 24394 48124 24400 48136
rect 24075 48096 24400 48124
rect 24075 48093 24087 48096
rect 24029 48087 24087 48093
rect 24394 48084 24400 48096
rect 24452 48084 24458 48136
rect 25222 48084 25228 48136
rect 25280 48084 25286 48136
rect 10459 47991 10517 47997
rect 10459 47957 10471 47991
rect 10505 47988 10517 47991
rect 12618 47988 12624 48000
rect 10505 47960 12624 47988
rect 10505 47957 10517 47960
rect 10459 47951 10517 47957
rect 12618 47948 12624 47960
rect 12676 47948 12682 48000
rect 21818 47948 21824 48000
rect 21876 47988 21882 48000
rect 23385 47991 23443 47997
rect 23385 47988 23397 47991
rect 21876 47960 23397 47988
rect 21876 47948 21882 47960
rect 23385 47957 23397 47960
rect 23431 47957 23443 47991
rect 23385 47951 23443 47957
rect 25133 47991 25191 47997
rect 25133 47957 25145 47991
rect 25179 47988 25191 47991
rect 25866 47988 25872 48000
rect 25179 47960 25872 47988
rect 25179 47957 25191 47960
rect 25133 47951 25191 47957
rect 25866 47948 25872 47960
rect 25924 47948 25930 48000
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9398 47744 9404 47796
rect 9456 47784 9462 47796
rect 9861 47787 9919 47793
rect 9861 47784 9873 47787
rect 9456 47756 9873 47784
rect 9456 47744 9462 47756
rect 9861 47753 9873 47756
rect 9907 47753 9919 47787
rect 9861 47747 9919 47753
rect 8478 47676 8484 47728
rect 8536 47716 8542 47728
rect 10137 47719 10195 47725
rect 10137 47716 10149 47719
rect 8536 47688 10149 47716
rect 8536 47676 8542 47688
rect 9416 47657 9444 47688
rect 10137 47685 10149 47688
rect 10183 47716 10195 47719
rect 10778 47716 10784 47728
rect 10183 47688 10784 47716
rect 10183 47685 10195 47688
rect 10137 47679 10195 47685
rect 10778 47676 10784 47688
rect 10836 47676 10842 47728
rect 9401 47651 9459 47657
rect 9401 47617 9413 47651
rect 9447 47648 9459 47651
rect 24857 47651 24915 47657
rect 9447 47620 9481 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 24857 47617 24869 47651
rect 24903 47648 24915 47651
rect 25314 47648 25320 47660
rect 24903 47620 25320 47648
rect 24903 47617 24915 47620
rect 24857 47611 24915 47617
rect 25314 47608 25320 47620
rect 25372 47608 25378 47660
rect 8846 47404 8852 47456
rect 8904 47444 8910 47456
rect 9122 47444 9128 47456
rect 8904 47416 9128 47444
rect 8904 47404 8910 47416
rect 9122 47404 9128 47416
rect 9180 47444 9186 47456
rect 9493 47447 9551 47453
rect 9493 47444 9505 47447
rect 9180 47416 9505 47444
rect 9180 47404 9186 47416
rect 9493 47413 9505 47416
rect 9539 47413 9551 47447
rect 9493 47407 9551 47413
rect 25133 47447 25191 47453
rect 25133 47413 25145 47447
rect 25179 47444 25191 47447
rect 25406 47444 25412 47456
rect 25179 47416 25412 47444
rect 25179 47413 25191 47416
rect 25133 47407 25191 47413
rect 25406 47404 25412 47416
rect 25464 47404 25470 47456
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 9398 46996 9404 47048
rect 9456 47036 9462 47048
rect 11644 47039 11702 47045
rect 11644 47036 11656 47039
rect 9456 47008 11656 47036
rect 9456 46996 9462 47008
rect 11644 47005 11656 47008
rect 11690 47005 11702 47039
rect 11644 46999 11702 47005
rect 11747 46971 11805 46977
rect 11747 46937 11759 46971
rect 11793 46968 11805 46971
rect 13722 46968 13728 46980
rect 11793 46940 13728 46968
rect 11793 46937 11805 46940
rect 11747 46931 11805 46937
rect 13722 46928 13728 46940
rect 13780 46928 13786 46980
rect 25314 46860 25320 46912
rect 25372 46900 25378 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 25372 46872 25421 46900
rect 25372 46860 25378 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 9766 46656 9772 46708
rect 9824 46696 9830 46708
rect 10318 46696 10324 46708
rect 9824 46668 10324 46696
rect 9824 46656 9830 46668
rect 10318 46656 10324 46668
rect 10376 46656 10382 46708
rect 10778 46656 10784 46708
rect 10836 46696 10842 46708
rect 11054 46696 11060 46708
rect 10836 46668 11060 46696
rect 10836 46656 10842 46668
rect 11054 46656 11060 46668
rect 11112 46656 11118 46708
rect 10336 46628 10364 46656
rect 10336 46600 11008 46628
rect 10778 46520 10784 46572
rect 10836 46520 10842 46572
rect 10980 46560 11008 46600
rect 13722 46588 13728 46640
rect 13780 46628 13786 46640
rect 14093 46631 14151 46637
rect 14093 46628 14105 46631
rect 13780 46600 14105 46628
rect 13780 46588 13786 46600
rect 14093 46597 14105 46600
rect 14139 46597 14151 46631
rect 14093 46591 14151 46597
rect 12564 46563 12622 46569
rect 12564 46560 12576 46563
rect 10980 46532 12576 46560
rect 12564 46529 12576 46532
rect 12610 46529 12622 46563
rect 12564 46523 12622 46529
rect 13906 46520 13912 46572
rect 13964 46520 13970 46572
rect 25314 46520 25320 46572
rect 25372 46520 25378 46572
rect 15746 46452 15752 46504
rect 15804 46452 15810 46504
rect 10594 46316 10600 46368
rect 10652 46316 10658 46368
rect 12667 46359 12725 46365
rect 12667 46325 12679 46359
rect 12713 46356 12725 46359
rect 16482 46356 16488 46368
rect 12713 46328 16488 46356
rect 12713 46325 12725 46328
rect 12667 46319 12725 46325
rect 16482 46316 16488 46328
rect 16540 46316 16546 46368
rect 25038 46316 25044 46368
rect 25096 46356 25102 46368
rect 25133 46359 25191 46365
rect 25133 46356 25145 46359
rect 25096 46328 25145 46356
rect 25096 46316 25102 46328
rect 25133 46325 25145 46328
rect 25179 46325 25191 46359
rect 25133 46319 25191 46325
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 7834 46112 7840 46164
rect 7892 46152 7898 46164
rect 7929 46155 7987 46161
rect 7929 46152 7941 46155
rect 7892 46124 7941 46152
rect 7892 46112 7898 46124
rect 7929 46121 7941 46124
rect 7975 46121 7987 46155
rect 7929 46115 7987 46121
rect 21726 46084 21732 46096
rect 16546 46056 21732 46084
rect 8389 46019 8447 46025
rect 8389 45985 8401 46019
rect 8435 46016 8447 46019
rect 9490 46016 9496 46028
rect 8435 45988 9496 46016
rect 8435 45985 8447 45988
rect 8389 45979 8447 45985
rect 9490 45976 9496 45988
rect 9548 45976 9554 46028
rect 16209 46019 16267 46025
rect 16209 45985 16221 46019
rect 16255 46016 16267 46019
rect 16546 46016 16574 46056
rect 21726 46044 21732 46056
rect 21784 46044 21790 46096
rect 16255 45988 16574 46016
rect 16669 46019 16727 46025
rect 16255 45985 16267 45988
rect 16209 45979 16267 45985
rect 16669 45985 16681 46019
rect 16715 46016 16727 46019
rect 16850 46016 16856 46028
rect 16715 45988 16856 46016
rect 16715 45985 16727 45988
rect 16669 45979 16727 45985
rect 16850 45976 16856 45988
rect 16908 45976 16914 46028
rect 8570 45908 8576 45960
rect 8628 45908 8634 45960
rect 10410 45908 10416 45960
rect 10468 45948 10474 45960
rect 13300 45951 13358 45957
rect 13300 45948 13312 45951
rect 10468 45920 13312 45948
rect 10468 45908 10474 45920
rect 13300 45917 13312 45920
rect 13346 45917 13358 45951
rect 13300 45911 13358 45917
rect 24857 45951 24915 45957
rect 24857 45917 24869 45951
rect 24903 45948 24915 45951
rect 25314 45948 25320 45960
rect 24903 45920 25320 45948
rect 24903 45917 24915 45920
rect 24857 45911 24915 45917
rect 25314 45908 25320 45920
rect 25372 45908 25378 45960
rect 16482 45840 16488 45892
rect 16540 45840 16546 45892
rect 13403 45815 13461 45821
rect 13403 45781 13415 45815
rect 13449 45812 13461 45815
rect 15102 45812 15108 45824
rect 13449 45784 15108 45812
rect 13449 45781 13461 45784
rect 13403 45775 13461 45781
rect 15102 45772 15108 45784
rect 15160 45772 15166 45824
rect 24946 45772 24952 45824
rect 25004 45812 25010 45824
rect 25133 45815 25191 45821
rect 25133 45812 25145 45815
rect 25004 45784 25145 45812
rect 25004 45772 25010 45784
rect 25133 45781 25145 45784
rect 25179 45781 25191 45815
rect 25133 45775 25191 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 12618 45500 12624 45552
rect 12676 45540 12682 45552
rect 12897 45543 12955 45549
rect 12897 45540 12909 45543
rect 12676 45512 12909 45540
rect 12676 45500 12682 45512
rect 12897 45509 12909 45512
rect 12943 45509 12955 45543
rect 12897 45503 12955 45509
rect 12710 45432 12716 45484
rect 12768 45432 12774 45484
rect 14550 45364 14556 45416
rect 14608 45364 14614 45416
rect 25314 45228 25320 45280
rect 25372 45268 25378 45280
rect 25409 45271 25467 45277
rect 25409 45268 25421 45271
rect 25372 45240 25421 45268
rect 25372 45228 25378 45240
rect 25409 45237 25421 45240
rect 25455 45237 25467 45271
rect 25409 45231 25467 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 9122 45024 9128 45076
rect 9180 45024 9186 45076
rect 19978 44996 19984 45008
rect 17052 44968 19984 44996
rect 17052 44937 17080 44968
rect 19978 44956 19984 44968
rect 20036 44956 20042 45008
rect 17037 44931 17095 44937
rect 17037 44897 17049 44931
rect 17083 44897 17095 44931
rect 17037 44891 17095 44897
rect 17494 44888 17500 44940
rect 17552 44888 17558 44940
rect 10870 44820 10876 44872
rect 10928 44860 10934 44872
rect 10928 44832 11376 44860
rect 10928 44820 10934 44832
rect 10166 44764 10364 44792
rect 8662 44684 8668 44736
rect 8720 44724 8726 44736
rect 10336 44724 10364 44764
rect 10594 44752 10600 44804
rect 10652 44752 10658 44804
rect 11348 44736 11376 44832
rect 25314 44820 25320 44872
rect 25372 44820 25378 44872
rect 15102 44752 15108 44804
rect 15160 44792 15166 44804
rect 17313 44795 17371 44801
rect 17313 44792 17325 44795
rect 15160 44764 17325 44792
rect 15160 44752 15166 44764
rect 17313 44761 17325 44764
rect 17359 44761 17371 44795
rect 17313 44755 17371 44761
rect 11146 44724 11152 44736
rect 8720 44696 11152 44724
rect 8720 44684 8726 44696
rect 11146 44684 11152 44696
rect 11204 44684 11210 44736
rect 11330 44684 11336 44736
rect 11388 44684 11394 44736
rect 25133 44727 25191 44733
rect 25133 44693 25145 44727
rect 25179 44724 25191 44727
rect 25314 44724 25320 44736
rect 25179 44696 25320 44724
rect 25179 44693 25191 44696
rect 25133 44687 25191 44693
rect 25314 44684 25320 44696
rect 25372 44684 25378 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 9582 44480 9588 44532
rect 9640 44480 9646 44532
rect 9125 44387 9183 44393
rect 9125 44353 9137 44387
rect 9171 44384 9183 44387
rect 9214 44384 9220 44396
rect 9171 44356 9220 44384
rect 9171 44353 9183 44356
rect 9125 44347 9183 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 11054 44344 11060 44396
rect 11112 44384 11118 44396
rect 11517 44387 11575 44393
rect 11517 44384 11529 44387
rect 11112 44356 11529 44384
rect 11112 44344 11118 44356
rect 11517 44353 11529 44356
rect 11563 44353 11575 44387
rect 11517 44347 11575 44353
rect 24765 44387 24823 44393
rect 24765 44353 24777 44387
rect 24811 44384 24823 44387
rect 25222 44384 25228 44396
rect 24811 44356 25228 44384
rect 24811 44353 24823 44356
rect 24765 44347 24823 44353
rect 25222 44344 25228 44356
rect 25280 44344 25286 44396
rect 8938 44276 8944 44328
rect 8996 44276 9002 44328
rect 10410 44140 10416 44192
rect 10468 44180 10474 44192
rect 10597 44183 10655 44189
rect 10597 44180 10609 44183
rect 10468 44152 10609 44180
rect 10468 44140 10474 44152
rect 10597 44149 10609 44152
rect 10643 44149 10655 44183
rect 10597 44143 10655 44149
rect 10962 44140 10968 44192
rect 11020 44140 11026 44192
rect 25133 44183 25191 44189
rect 25133 44149 25145 44183
rect 25179 44180 25191 44183
rect 25682 44180 25688 44192
rect 25179 44152 25688 44180
rect 25179 44149 25191 44152
rect 25133 44143 25191 44149
rect 25682 44140 25688 44152
rect 25740 44140 25746 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 21818 43800 21824 43852
rect 21876 43800 21882 43852
rect 20714 43732 20720 43784
rect 20772 43732 20778 43784
rect 22097 43775 22155 43781
rect 22097 43741 22109 43775
rect 22143 43772 22155 43775
rect 23382 43772 23388 43784
rect 22143 43744 23388 43772
rect 22143 43741 22155 43744
rect 22097 43735 22155 43741
rect 23382 43732 23388 43744
rect 23440 43732 23446 43784
rect 16574 43596 16580 43648
rect 16632 43636 16638 43648
rect 20349 43639 20407 43645
rect 20349 43636 20361 43639
rect 16632 43608 20361 43636
rect 16632 43596 16638 43608
rect 20349 43605 20361 43608
rect 20395 43605 20407 43639
rect 20732 43636 20760 43732
rect 22373 43639 22431 43645
rect 22373 43636 22385 43639
rect 20732 43608 22385 43636
rect 20349 43599 20407 43605
rect 22373 43605 22385 43608
rect 22419 43605 22431 43639
rect 22373 43599 22431 43605
rect 25222 43596 25228 43648
rect 25280 43636 25286 43648
rect 25409 43639 25467 43645
rect 25409 43636 25421 43639
rect 25280 43608 25421 43636
rect 25280 43596 25286 43608
rect 25409 43605 25421 43608
rect 25455 43605 25467 43639
rect 25409 43599 25467 43605
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 25222 43256 25228 43308
rect 25280 43256 25286 43308
rect 24302 43120 24308 43172
rect 24360 43160 24366 43172
rect 25041 43163 25099 43169
rect 25041 43160 25053 43163
rect 24360 43132 25053 43160
rect 24360 43120 24366 43132
rect 25041 43129 25053 43132
rect 25087 43129 25099 43163
rect 25041 43123 25099 43129
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 9766 42712 9772 42764
rect 9824 42712 9830 42764
rect 10226 42712 10232 42764
rect 10284 42712 10290 42764
rect 9030 42644 9036 42696
rect 9088 42684 9094 42696
rect 9585 42687 9643 42693
rect 9585 42684 9597 42687
rect 9088 42656 9597 42684
rect 9088 42644 9094 42656
rect 9585 42653 9597 42656
rect 9631 42653 9643 42687
rect 9585 42647 9643 42653
rect 24765 42619 24823 42625
rect 24765 42585 24777 42619
rect 24811 42616 24823 42619
rect 25222 42616 25228 42628
rect 24811 42588 25228 42616
rect 24811 42585 24823 42588
rect 24765 42579 24823 42585
rect 25222 42576 25228 42588
rect 25280 42576 25286 42628
rect 20990 42508 20996 42560
rect 21048 42548 21054 42560
rect 25133 42551 25191 42557
rect 25133 42548 25145 42551
rect 21048 42520 25145 42548
rect 21048 42508 21054 42520
rect 25133 42517 25145 42520
rect 25179 42517 25191 42551
rect 25133 42511 25191 42517
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 9401 42347 9459 42353
rect 9401 42313 9413 42347
rect 9447 42344 9459 42347
rect 10594 42344 10600 42356
rect 9447 42316 10600 42344
rect 9447 42313 9459 42316
rect 9401 42307 9459 42313
rect 10594 42304 10600 42316
rect 10652 42304 10658 42356
rect 11146 42344 11152 42356
rect 10704 42316 11152 42344
rect 10704 42276 10732 42316
rect 11146 42304 11152 42316
rect 11204 42344 11210 42356
rect 11514 42344 11520 42356
rect 11204 42316 11520 42344
rect 11204 42304 11210 42316
rect 11514 42304 11520 42316
rect 11572 42304 11578 42356
rect 10442 42248 10732 42276
rect 10873 42279 10931 42285
rect 10873 42245 10885 42279
rect 10919 42276 10931 42279
rect 10962 42276 10968 42288
rect 10919 42248 10968 42276
rect 10919 42245 10931 42248
rect 10873 42239 10931 42245
rect 10962 42236 10968 42248
rect 11020 42236 11026 42288
rect 11149 42143 11207 42149
rect 11149 42109 11161 42143
rect 11195 42140 11207 42143
rect 11330 42140 11336 42152
rect 11195 42112 11336 42140
rect 11195 42109 11207 42112
rect 11149 42103 11207 42109
rect 11330 42100 11336 42112
rect 11388 42140 11394 42152
rect 11388 42112 11744 42140
rect 11388 42100 11394 42112
rect 11716 42016 11744 42112
rect 11514 41964 11520 42016
rect 11572 41964 11578 42016
rect 11698 41964 11704 42016
rect 11756 41964 11762 42016
rect 25222 41964 25228 42016
rect 25280 42004 25286 42016
rect 25409 42007 25467 42013
rect 25409 42004 25421 42007
rect 25280 41976 25421 42004
rect 25280 41964 25286 41976
rect 25409 41973 25421 41976
rect 25455 41973 25467 42007
rect 25409 41967 25467 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 10870 41760 10876 41812
rect 10928 41760 10934 41812
rect 10410 41624 10416 41676
rect 10468 41624 10474 41676
rect 10226 41556 10232 41608
rect 10284 41556 10290 41608
rect 25222 41556 25228 41608
rect 25280 41556 25286 41608
rect 24854 41488 24860 41540
rect 24912 41528 24918 41540
rect 25041 41531 25099 41537
rect 25041 41528 25053 41531
rect 24912 41500 25053 41528
rect 24912 41488 24918 41500
rect 25041 41497 25053 41500
rect 25087 41497 25099 41531
rect 25041 41491 25099 41497
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 24857 41123 24915 41129
rect 24857 41089 24869 41123
rect 24903 41120 24915 41123
rect 25314 41120 25320 41132
rect 24903 41092 25320 41120
rect 24903 41089 24915 41092
rect 24857 41083 24915 41089
rect 25314 41080 25320 41092
rect 25372 41080 25378 41132
rect 24854 40876 24860 40928
rect 24912 40916 24918 40928
rect 25038 40916 25044 40928
rect 24912 40888 25044 40916
rect 24912 40876 24918 40888
rect 25038 40876 25044 40888
rect 25096 40876 25102 40928
rect 25133 40919 25191 40925
rect 25133 40885 25145 40919
rect 25179 40916 25191 40919
rect 26602 40916 26608 40928
rect 25179 40888 26608 40916
rect 25179 40885 25191 40888
rect 25133 40879 25191 40885
rect 26602 40876 26608 40888
rect 26660 40876 26666 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 24946 40332 24952 40384
rect 25004 40372 25010 40384
rect 25222 40372 25228 40384
rect 25004 40344 25228 40372
rect 25004 40332 25010 40344
rect 25222 40332 25228 40344
rect 25280 40332 25286 40384
rect 25498 40332 25504 40384
rect 25556 40332 25562 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 23290 40128 23296 40180
rect 23348 40168 23354 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 23348 40140 25145 40168
rect 23348 40128 23354 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 25498 40100 25504 40112
rect 25332 40072 25504 40100
rect 25332 40041 25360 40072
rect 25498 40060 25504 40072
rect 25556 40060 25562 40112
rect 25317 40035 25375 40041
rect 25317 40001 25329 40035
rect 25363 40001 25375 40035
rect 25317 39995 25375 40001
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39420 24915 39423
rect 25314 39420 25320 39432
rect 24903 39392 25320 39420
rect 24903 39389 24915 39392
rect 24857 39383 24915 39389
rect 25314 39380 25320 39392
rect 25372 39380 25378 39432
rect 22002 39244 22008 39296
rect 22060 39284 22066 39296
rect 25133 39287 25191 39293
rect 25133 39284 25145 39287
rect 22060 39256 25145 39284
rect 22060 39244 22066 39256
rect 25133 39253 25145 39256
rect 25179 39253 25191 39287
rect 25133 39247 25191 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25409 38743 25467 38749
rect 25409 38740 25421 38743
rect 25372 38712 25421 38740
rect 25372 38700 25378 38712
rect 25409 38709 25421 38712
rect 25455 38709 25467 38743
rect 25409 38703 25467 38709
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 25314 38292 25320 38344
rect 25372 38292 25378 38344
rect 25133 38199 25191 38205
rect 25133 38165 25145 38199
rect 25179 38196 25191 38199
rect 25498 38196 25504 38208
rect 25179 38168 25504 38196
rect 25179 38165 25191 38168
rect 25133 38159 25191 38165
rect 25498 38156 25504 38168
rect 25556 38156 25562 38208
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 8570 37952 8576 38004
rect 8628 37992 8634 38004
rect 8665 37995 8723 38001
rect 8665 37992 8677 37995
rect 8628 37964 8677 37992
rect 8628 37952 8634 37964
rect 8665 37961 8677 37964
rect 8711 37961 8723 37995
rect 8665 37955 8723 37961
rect 8846 37816 8852 37868
rect 8904 37816 8910 37868
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 25222 37856 25228 37868
rect 24811 37828 25228 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 25222 37816 25228 37828
rect 25280 37816 25286 37868
rect 25133 37655 25191 37661
rect 25133 37621 25145 37655
rect 25179 37652 25191 37655
rect 25958 37652 25964 37664
rect 25179 37624 25964 37652
rect 25179 37621 25191 37624
rect 25133 37615 25191 37621
rect 25958 37612 25964 37624
rect 26016 37612 26022 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 25222 37068 25228 37120
rect 25280 37108 25286 37120
rect 25409 37111 25467 37117
rect 25409 37108 25421 37111
rect 25280 37080 25421 37108
rect 25280 37068 25286 37080
rect 25409 37077 25421 37080
rect 25455 37077 25467 37111
rect 25409 37071 25467 37077
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 25222 36728 25228 36780
rect 25280 36728 25286 36780
rect 25133 36567 25191 36573
rect 25133 36533 25145 36567
rect 25179 36564 25191 36567
rect 25774 36564 25780 36576
rect 25179 36536 25780 36564
rect 25179 36533 25191 36536
rect 25133 36527 25191 36533
rect 25774 36524 25780 36536
rect 25832 36524 25838 36576
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 36020 25191 36023
rect 26786 36020 26792 36032
rect 25179 35992 26792 36020
rect 25179 35989 25191 35992
rect 25133 35983 25191 35989
rect 26786 35980 26792 35992
rect 26844 35980 26850 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 11698 35816 11704 35828
rect 9416 35788 11704 35816
rect 9416 35689 9444 35788
rect 11698 35776 11704 35788
rect 11756 35776 11762 35828
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 25038 35816 25044 35828
rect 22511 35788 25044 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 25038 35776 25044 35788
rect 25096 35776 25102 35828
rect 11514 35748 11520 35760
rect 10902 35720 11520 35748
rect 11514 35708 11520 35720
rect 11572 35708 11578 35760
rect 21177 35751 21235 35757
rect 21177 35717 21189 35751
rect 21223 35748 21235 35751
rect 24854 35748 24860 35760
rect 21223 35720 24860 35748
rect 21223 35717 21235 35720
rect 21177 35711 21235 35717
rect 24854 35708 24860 35720
rect 24912 35708 24918 35760
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35649 9459 35683
rect 9401 35643 9459 35649
rect 15746 35640 15752 35692
rect 15804 35680 15810 35692
rect 20441 35683 20499 35689
rect 20441 35680 20453 35683
rect 15804 35652 20453 35680
rect 15804 35640 15810 35652
rect 20441 35649 20453 35652
rect 20487 35680 20499 35683
rect 21082 35680 21088 35692
rect 20487 35652 21088 35680
rect 20487 35649 20499 35652
rect 20441 35643 20499 35649
rect 21082 35640 21088 35652
rect 21140 35640 21146 35692
rect 21726 35640 21732 35692
rect 21784 35680 21790 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 21784 35652 22385 35680
rect 21784 35640 21790 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 11149 35615 11207 35621
rect 11149 35612 11161 35615
rect 11020 35584 11161 35612
rect 11020 35572 11026 35584
rect 11149 35581 11161 35584
rect 11195 35581 11207 35615
rect 11149 35575 11207 35581
rect 21266 35572 21272 35624
rect 21324 35572 21330 35624
rect 22554 35572 22560 35624
rect 22612 35572 22618 35624
rect 19242 35504 19248 35556
rect 19300 35544 19306 35556
rect 19300 35516 20484 35544
rect 19300 35504 19306 35516
rect 11790 35436 11796 35488
rect 11848 35436 11854 35488
rect 20456 35476 20484 35516
rect 20530 35504 20536 35556
rect 20588 35544 20594 35556
rect 22005 35547 22063 35553
rect 22005 35544 22017 35547
rect 20588 35516 22017 35544
rect 20588 35504 20594 35516
rect 22005 35513 22017 35516
rect 22051 35513 22063 35547
rect 22005 35507 22063 35513
rect 20717 35479 20775 35485
rect 20717 35476 20729 35479
rect 20456 35448 20729 35476
rect 20717 35445 20729 35448
rect 20763 35445 20775 35479
rect 20717 35439 20775 35445
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 21726 35232 21732 35284
rect 21784 35272 21790 35284
rect 21821 35275 21879 35281
rect 21821 35272 21833 35275
rect 21784 35244 21833 35272
rect 21784 35232 21790 35244
rect 21821 35241 21833 35244
rect 21867 35241 21879 35275
rect 21821 35235 21879 35241
rect 22278 35096 22284 35148
rect 22336 35136 22342 35148
rect 23293 35139 23351 35145
rect 23293 35136 23305 35139
rect 22336 35108 23305 35136
rect 22336 35096 22342 35108
rect 23293 35105 23305 35108
rect 23339 35105 23351 35139
rect 23293 35099 23351 35105
rect 23201 35071 23259 35077
rect 23201 35037 23213 35071
rect 23247 35068 23259 35071
rect 24946 35068 24952 35080
rect 23247 35040 24952 35068
rect 23247 35037 23259 35040
rect 23201 35031 23259 35037
rect 24946 35028 24952 35040
rect 25004 35028 25010 35080
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 20254 35000 20260 35012
rect 20036 34972 20260 35000
rect 20036 34960 20042 34972
rect 20254 34960 20260 34972
rect 20312 35000 20318 35012
rect 22373 35003 22431 35009
rect 22373 35000 22385 35003
rect 20312 34972 22385 35000
rect 20312 34960 20318 34972
rect 22373 34969 22385 34972
rect 22419 35000 22431 35003
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 22419 34972 23121 35000
rect 22419 34969 22431 34972
rect 22373 34963 22431 34969
rect 23109 34969 23121 34972
rect 23155 34969 23167 35003
rect 23109 34963 23167 34969
rect 22738 34892 22744 34944
rect 22796 34892 22802 34944
rect 25133 34935 25191 34941
rect 25133 34901 25145 34935
rect 25179 34932 25191 34935
rect 26142 34932 26148 34944
rect 25179 34904 26148 34932
rect 25179 34901 25191 34904
rect 25133 34895 25191 34901
rect 26142 34892 26148 34904
rect 26200 34892 26206 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 20346 34688 20352 34740
rect 20404 34728 20410 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 20404 34700 25145 34728
rect 20404 34688 20410 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 24857 34595 24915 34601
rect 24857 34561 24869 34595
rect 24903 34592 24915 34595
rect 25314 34592 25320 34604
rect 24903 34564 25320 34592
rect 24903 34561 24915 34564
rect 24857 34555 24915 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 20714 34348 20720 34400
rect 20772 34388 20778 34400
rect 21361 34391 21419 34397
rect 21361 34388 21373 34391
rect 20772 34360 21373 34388
rect 20772 34348 20778 34360
rect 21361 34357 21373 34360
rect 21407 34388 21419 34391
rect 21818 34388 21824 34400
rect 21407 34360 21824 34388
rect 21407 34357 21419 34360
rect 21361 34351 21419 34357
rect 21818 34348 21824 34360
rect 21876 34348 21882 34400
rect 22186 34348 22192 34400
rect 22244 34388 22250 34400
rect 22646 34388 22652 34400
rect 22244 34360 22652 34388
rect 22244 34348 22250 34360
rect 22646 34348 22652 34360
rect 22704 34348 22710 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 8938 34144 8944 34196
rect 8996 34184 9002 34196
rect 9125 34187 9183 34193
rect 9125 34184 9137 34187
rect 8996 34156 9137 34184
rect 8996 34144 9002 34156
rect 9125 34153 9137 34156
rect 9171 34153 9183 34187
rect 9125 34147 9183 34153
rect 21637 34187 21695 34193
rect 21637 34153 21649 34187
rect 21683 34184 21695 34187
rect 22094 34184 22100 34196
rect 21683 34156 22100 34184
rect 21683 34153 21695 34156
rect 21637 34147 21695 34153
rect 22094 34144 22100 34156
rect 22152 34184 22158 34196
rect 22554 34184 22560 34196
rect 22152 34156 22560 34184
rect 22152 34144 22158 34156
rect 22554 34144 22560 34156
rect 22612 34144 22618 34196
rect 11790 34008 11796 34060
rect 11848 34048 11854 34060
rect 14737 34051 14795 34057
rect 14737 34048 14749 34051
rect 11848 34020 14749 34048
rect 11848 34008 11854 34020
rect 14737 34017 14749 34020
rect 14783 34017 14795 34051
rect 14737 34011 14795 34017
rect 22646 34008 22652 34060
rect 22704 34048 22710 34060
rect 23109 34051 23167 34057
rect 23109 34048 23121 34051
rect 22704 34020 23121 34048
rect 22704 34008 22710 34020
rect 23109 34017 23121 34020
rect 23155 34017 23167 34051
rect 23109 34011 23167 34017
rect 23382 34008 23388 34060
rect 23440 34008 23446 34060
rect 9214 33940 9220 33992
rect 9272 33980 9278 33992
rect 9309 33983 9367 33989
rect 9309 33980 9321 33983
rect 9272 33952 9321 33980
rect 9272 33940 9278 33952
rect 9309 33949 9321 33952
rect 9355 33949 9367 33983
rect 9309 33943 9367 33949
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 19429 33983 19487 33989
rect 19429 33980 19441 33983
rect 19392 33952 19441 33980
rect 19392 33940 19398 33952
rect 19429 33949 19441 33952
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 15565 33915 15623 33921
rect 15565 33881 15577 33915
rect 15611 33912 15623 33915
rect 15841 33915 15899 33921
rect 15841 33912 15853 33915
rect 15611 33884 15853 33912
rect 15611 33881 15623 33884
rect 15565 33875 15623 33881
rect 15841 33881 15853 33884
rect 15887 33912 15899 33915
rect 16298 33912 16304 33924
rect 15887 33884 16304 33912
rect 15887 33881 15899 33884
rect 15841 33875 15899 33881
rect 16298 33872 16304 33884
rect 16356 33872 16362 33924
rect 19702 33872 19708 33924
rect 19760 33872 19766 33924
rect 20162 33872 20168 33924
rect 20220 33872 20226 33924
rect 21818 33872 21824 33924
rect 21876 33912 21882 33924
rect 21876 33884 21942 33912
rect 21876 33872 21882 33884
rect 23198 33872 23204 33924
rect 23256 33912 23262 33924
rect 23400 33912 23428 34008
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25314 33980 25320 33992
rect 24903 33952 25320 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 23256 33884 23428 33912
rect 23256 33872 23262 33884
rect 21174 33804 21180 33856
rect 21232 33804 21238 33856
rect 23753 33847 23811 33853
rect 23753 33813 23765 33847
rect 23799 33844 23811 33847
rect 24210 33844 24216 33856
rect 23799 33816 24216 33844
rect 23799 33813 23811 33816
rect 23753 33807 23811 33813
rect 24210 33804 24216 33816
rect 24268 33804 24274 33856
rect 25133 33847 25191 33853
rect 25133 33813 25145 33847
rect 25179 33844 25191 33847
rect 26234 33844 26240 33856
rect 25179 33816 26240 33844
rect 25179 33813 25191 33816
rect 25133 33807 25191 33813
rect 26234 33804 26240 33816
rect 26292 33804 26298 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 20162 33600 20168 33652
rect 20220 33640 20226 33652
rect 21637 33643 21695 33649
rect 21637 33640 21649 33643
rect 20220 33612 21649 33640
rect 20220 33600 20226 33612
rect 20640 33572 20668 33612
rect 21637 33609 21649 33612
rect 21683 33640 21695 33643
rect 21818 33640 21824 33652
rect 21683 33612 21824 33640
rect 21683 33609 21695 33612
rect 21637 33603 21695 33609
rect 21818 33600 21824 33612
rect 21876 33640 21882 33652
rect 21876 33612 22416 33640
rect 21876 33600 21882 33612
rect 20562 33544 20668 33572
rect 22278 33532 22284 33584
rect 22336 33532 22342 33584
rect 22388 33572 22416 33612
rect 22554 33600 22560 33652
rect 22612 33640 22618 33652
rect 23753 33643 23811 33649
rect 23753 33640 23765 33643
rect 22612 33612 23765 33640
rect 22612 33600 22618 33612
rect 23753 33609 23765 33612
rect 23799 33609 23811 33643
rect 23753 33603 23811 33609
rect 22388 33544 22770 33572
rect 25317 33507 25375 33513
rect 25317 33504 25329 33507
rect 24872 33476 25329 33504
rect 20993 33439 21051 33445
rect 20993 33405 21005 33439
rect 21039 33436 21051 33439
rect 21269 33439 21327 33445
rect 21039 33408 21220 33436
rect 21039 33405 21051 33408
rect 20993 33399 21051 33405
rect 19521 33303 19579 33309
rect 19521 33269 19533 33303
rect 19567 33300 19579 33303
rect 19702 33300 19708 33312
rect 19567 33272 19708 33300
rect 19567 33269 19579 33272
rect 19521 33263 19579 33269
rect 19702 33260 19708 33272
rect 19760 33300 19766 33312
rect 20438 33300 20444 33312
rect 19760 33272 20444 33300
rect 19760 33260 19766 33272
rect 20438 33260 20444 33272
rect 20496 33260 20502 33312
rect 21192 33300 21220 33408
rect 21269 33405 21281 33439
rect 21315 33436 21327 33439
rect 22005 33439 22063 33445
rect 22005 33436 22017 33439
rect 21315 33408 22017 33436
rect 21315 33405 21327 33408
rect 21269 33399 21327 33405
rect 22005 33405 22017 33408
rect 22051 33436 22063 33439
rect 23290 33436 23296 33448
rect 22051 33408 23296 33436
rect 22051 33405 22063 33408
rect 22005 33399 22063 33405
rect 23290 33396 23296 33408
rect 23348 33396 23354 33448
rect 22094 33300 22100 33312
rect 21192 33272 22100 33300
rect 22094 33260 22100 33272
rect 22152 33260 22158 33312
rect 24210 33260 24216 33312
rect 24268 33300 24274 33312
rect 24305 33303 24363 33309
rect 24305 33300 24317 33303
rect 24268 33272 24317 33300
rect 24268 33260 24274 33272
rect 24305 33269 24317 33272
rect 24351 33269 24363 33303
rect 24305 33263 24363 33269
rect 24578 33260 24584 33312
rect 24636 33260 24642 33312
rect 24762 33260 24768 33312
rect 24820 33300 24826 33312
rect 24872 33309 24900 33476
rect 25317 33473 25329 33476
rect 25363 33473 25375 33507
rect 25317 33467 25375 33473
rect 25406 33328 25412 33380
rect 25464 33368 25470 33380
rect 26418 33368 26424 33380
rect 25464 33340 26424 33368
rect 25464 33328 25470 33340
rect 26418 33328 26424 33340
rect 26476 33328 26482 33380
rect 24857 33303 24915 33309
rect 24857 33300 24869 33303
rect 24820 33272 24869 33300
rect 24820 33260 24826 33272
rect 24857 33269 24869 33272
rect 24903 33269 24915 33303
rect 24857 33263 24915 33269
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 26050 33300 26056 33312
rect 25179 33272 26056 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 26050 33260 26056 33272
rect 26108 33260 26114 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 16758 33056 16764 33108
rect 16816 33096 16822 33108
rect 17310 33096 17316 33108
rect 16816 33068 17316 33096
rect 16816 33056 16822 33068
rect 17310 33056 17316 33068
rect 17368 33056 17374 33108
rect 22278 33056 22284 33108
rect 22336 33056 22342 33108
rect 23566 33096 23572 33108
rect 22388 33068 23572 33096
rect 17037 33031 17095 33037
rect 17037 32997 17049 33031
rect 17083 33028 17095 33031
rect 22388 33028 22416 33068
rect 23566 33056 23572 33068
rect 23624 33056 23630 33108
rect 17083 33000 22416 33028
rect 17083 32997 17095 33000
rect 17037 32991 17095 32997
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 16574 32960 16580 32972
rect 16264 32932 16580 32960
rect 16264 32920 16270 32932
rect 16574 32920 16580 32932
rect 16632 32960 16638 32972
rect 16632 32932 16677 32960
rect 16632 32920 16638 32932
rect 16025 32895 16083 32901
rect 16025 32861 16037 32895
rect 16071 32892 16083 32895
rect 16758 32892 16764 32904
rect 16071 32864 16764 32892
rect 16071 32861 16083 32864
rect 16025 32855 16083 32861
rect 16758 32852 16764 32864
rect 16816 32852 16822 32904
rect 15933 32827 15991 32833
rect 15933 32793 15945 32827
rect 15979 32824 15991 32827
rect 15979 32796 16574 32824
rect 15979 32793 15991 32796
rect 15933 32787 15991 32793
rect 12618 32716 12624 32768
rect 12676 32756 12682 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 12676 32728 15577 32756
rect 12676 32716 12682 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 16546 32756 16574 32796
rect 17052 32756 17080 32991
rect 23290 32920 23296 32972
rect 23348 32960 23354 32972
rect 24029 32963 24087 32969
rect 24029 32960 24041 32963
rect 23348 32932 24041 32960
rect 23348 32920 23354 32932
rect 24029 32929 24041 32932
rect 24075 32929 24087 32963
rect 24029 32923 24087 32929
rect 24765 32963 24823 32969
rect 24765 32929 24777 32963
rect 24811 32960 24823 32963
rect 24946 32960 24952 32972
rect 24811 32932 24952 32960
rect 24811 32929 24823 32932
rect 24765 32923 24823 32929
rect 24946 32920 24952 32932
rect 25004 32920 25010 32972
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 26602 32892 26608 32904
rect 24903 32864 26608 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 26602 32852 26608 32864
rect 26660 32852 26666 32904
rect 19889 32827 19947 32833
rect 19889 32793 19901 32827
rect 19935 32824 19947 32827
rect 20717 32827 20775 32833
rect 19935 32796 19969 32824
rect 19935 32793 19947 32796
rect 19889 32787 19947 32793
rect 20717 32793 20729 32827
rect 20763 32824 20775 32827
rect 20806 32824 20812 32836
rect 20763 32796 20812 32824
rect 20763 32793 20775 32796
rect 20717 32787 20775 32793
rect 17218 32756 17224 32768
rect 16546 32728 17224 32756
rect 15565 32719 15623 32725
rect 17218 32716 17224 32728
rect 17276 32716 17282 32768
rect 19613 32759 19671 32765
rect 19613 32725 19625 32759
rect 19659 32756 19671 32759
rect 19904 32756 19932 32787
rect 20806 32784 20812 32796
rect 20864 32784 20870 32836
rect 23198 32784 23204 32836
rect 23256 32784 23262 32836
rect 23753 32827 23811 32833
rect 23753 32793 23765 32827
rect 23799 32824 23811 32827
rect 25406 32824 25412 32836
rect 23799 32796 25412 32824
rect 23799 32793 23811 32796
rect 23753 32787 23811 32793
rect 25406 32784 25412 32796
rect 25464 32784 25470 32836
rect 21818 32756 21824 32768
rect 19659 32728 21824 32756
rect 19659 32725 19671 32728
rect 19613 32719 19671 32725
rect 21818 32716 21824 32728
rect 21876 32716 21882 32768
rect 24578 32716 24584 32768
rect 24636 32756 24642 32768
rect 24949 32759 25007 32765
rect 24949 32756 24961 32759
rect 24636 32728 24961 32756
rect 24636 32716 24642 32728
rect 24949 32725 24961 32728
rect 24995 32725 25007 32759
rect 24949 32719 25007 32725
rect 25222 32716 25228 32768
rect 25280 32756 25286 32768
rect 25317 32759 25375 32765
rect 25317 32756 25329 32759
rect 25280 32728 25329 32756
rect 25280 32716 25286 32728
rect 25317 32725 25329 32728
rect 25363 32725 25375 32759
rect 25317 32719 25375 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 16666 32512 16672 32564
rect 16724 32552 16730 32564
rect 16853 32555 16911 32561
rect 16853 32552 16865 32555
rect 16724 32524 16865 32552
rect 16724 32512 16730 32524
rect 16853 32521 16865 32524
rect 16899 32552 16911 32555
rect 23842 32552 23848 32564
rect 16899 32524 23848 32552
rect 16899 32521 16911 32524
rect 16853 32515 16911 32521
rect 23842 32512 23848 32524
rect 23900 32512 23906 32564
rect 16298 32444 16304 32496
rect 16356 32484 16362 32496
rect 16356 32456 16574 32484
rect 16356 32444 16362 32456
rect 16546 32416 16574 32456
rect 20070 32444 20076 32496
rect 20128 32444 20134 32496
rect 20533 32487 20591 32493
rect 20533 32453 20545 32487
rect 20579 32484 20591 32487
rect 21174 32484 21180 32496
rect 20579 32456 21180 32484
rect 20579 32453 20591 32456
rect 20533 32447 20591 32453
rect 21174 32444 21180 32456
rect 21232 32444 21238 32496
rect 23198 32444 23204 32496
rect 23256 32484 23262 32496
rect 23750 32484 23756 32496
rect 23256 32456 23756 32484
rect 23256 32444 23262 32456
rect 23750 32444 23756 32456
rect 23808 32484 23814 32496
rect 24210 32484 24216 32496
rect 23808 32456 24216 32484
rect 23808 32444 23814 32456
rect 24210 32444 24216 32456
rect 24268 32444 24274 32496
rect 16546 32388 17080 32416
rect 15470 32308 15476 32360
rect 15528 32308 15534 32360
rect 17052 32224 17080 32388
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 21876 32388 22109 32416
rect 21876 32376 21882 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 22462 32376 22468 32428
rect 22520 32416 22526 32428
rect 22925 32419 22983 32425
rect 22925 32416 22937 32419
rect 22520 32388 22937 32416
rect 22520 32376 22526 32388
rect 22925 32385 22937 32388
rect 22971 32416 22983 32419
rect 23290 32416 23296 32428
rect 22971 32388 23296 32416
rect 22971 32385 22983 32388
rect 22925 32379 22983 32385
rect 23290 32376 23296 32388
rect 23348 32416 23354 32428
rect 23477 32419 23535 32425
rect 23477 32416 23489 32419
rect 23348 32388 23489 32416
rect 23348 32376 23354 32388
rect 23477 32385 23489 32388
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 20806 32348 20812 32360
rect 20732 32320 20812 32348
rect 17034 32172 17040 32224
rect 17092 32172 17098 32224
rect 19058 32172 19064 32224
rect 19116 32172 19122 32224
rect 19426 32172 19432 32224
rect 19484 32212 19490 32224
rect 20732 32212 20760 32320
rect 20806 32308 20812 32320
rect 20864 32308 20870 32360
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 24946 32348 24952 32360
rect 23799 32320 24952 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 24946 32308 24952 32320
rect 25004 32308 25010 32360
rect 19484 32184 20760 32212
rect 19484 32172 19490 32184
rect 21082 32172 21088 32224
rect 21140 32172 21146 32224
rect 21637 32215 21695 32221
rect 21637 32181 21649 32215
rect 21683 32212 21695 32215
rect 21818 32212 21824 32224
rect 21683 32184 21824 32212
rect 21683 32181 21695 32184
rect 21637 32175 21695 32181
rect 21818 32172 21824 32184
rect 21876 32172 21882 32224
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 22830 32212 22836 32224
rect 22152 32184 22836 32212
rect 22152 32172 22158 32184
rect 22830 32172 22836 32184
rect 22888 32172 22894 32224
rect 25225 32215 25283 32221
rect 25225 32181 25237 32215
rect 25271 32212 25283 32215
rect 25406 32212 25412 32224
rect 25271 32184 25412 32212
rect 25271 32181 25283 32184
rect 25225 32175 25283 32181
rect 25406 32172 25412 32184
rect 25464 32172 25470 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 16850 31968 16856 32020
rect 16908 32008 16914 32020
rect 17402 32008 17408 32020
rect 16908 31980 17408 32008
rect 16908 31968 16914 31980
rect 17402 31968 17408 31980
rect 17460 31968 17466 32020
rect 20162 31968 20168 32020
rect 20220 32008 20226 32020
rect 21082 32008 21088 32020
rect 20220 31980 21088 32008
rect 20220 31968 20226 31980
rect 21082 31968 21088 31980
rect 21140 31968 21146 32020
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 15565 31943 15623 31949
rect 15565 31940 15577 31943
rect 12584 31912 15577 31940
rect 12584 31900 12590 31912
rect 15565 31909 15577 31912
rect 15611 31909 15623 31943
rect 16868 31940 16896 31968
rect 15565 31903 15623 31909
rect 16040 31912 16896 31940
rect 20732 31912 22232 31940
rect 16040 31881 16068 31912
rect 16025 31875 16083 31881
rect 16025 31841 16037 31875
rect 16071 31841 16083 31875
rect 16025 31835 16083 31841
rect 16206 31832 16212 31884
rect 16264 31832 16270 31884
rect 17770 31832 17776 31884
rect 17828 31872 17834 31884
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 17828 31844 18521 31872
rect 17828 31832 17834 31844
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 18509 31835 18567 31841
rect 19702 31832 19708 31884
rect 19760 31872 19766 31884
rect 20732 31872 20760 31912
rect 19760 31844 20760 31872
rect 19760 31832 19766 31844
rect 20898 31832 20904 31884
rect 20956 31872 20962 31884
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 20956 31844 21189 31872
rect 20956 31832 20962 31844
rect 21177 31841 21189 31844
rect 21223 31841 21235 31875
rect 21177 31835 21235 31841
rect 22002 31832 22008 31884
rect 22060 31872 22066 31884
rect 22204 31881 22232 31912
rect 22830 31900 22836 31952
rect 22888 31940 22894 31952
rect 23017 31943 23075 31949
rect 23017 31940 23029 31943
rect 22888 31912 23029 31940
rect 22888 31900 22894 31912
rect 23017 31909 23029 31912
rect 23063 31909 23075 31943
rect 23017 31903 23075 31909
rect 25038 31900 25044 31952
rect 25096 31940 25102 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 25096 31912 25145 31940
rect 25096 31900 25102 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 22097 31875 22155 31881
rect 22097 31872 22109 31875
rect 22060 31844 22109 31872
rect 22060 31832 22066 31844
rect 22097 31841 22109 31844
rect 22143 31841 22155 31875
rect 22097 31835 22155 31841
rect 22189 31875 22247 31881
rect 22189 31841 22201 31875
rect 22235 31841 22247 31875
rect 22189 31835 22247 31841
rect 23382 31832 23388 31884
rect 23440 31872 23446 31884
rect 23477 31875 23535 31881
rect 23477 31872 23489 31875
rect 23440 31844 23489 31872
rect 23440 31832 23446 31844
rect 23477 31841 23489 31844
rect 23523 31841 23535 31875
rect 23477 31835 23535 31841
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31841 23627 31875
rect 23569 31835 23627 31841
rect 15470 31764 15476 31816
rect 15528 31804 15534 31816
rect 16758 31804 16764 31816
rect 15528 31776 16764 31804
rect 15528 31764 15534 31776
rect 16758 31764 16764 31776
rect 16816 31764 16822 31816
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 23014 31764 23020 31816
rect 23072 31804 23078 31816
rect 23584 31804 23612 31835
rect 23072 31776 23612 31804
rect 24857 31807 24915 31813
rect 23072 31764 23078 31776
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 17037 31739 17095 31745
rect 17037 31705 17049 31739
rect 17083 31736 17095 31739
rect 17126 31736 17132 31748
rect 17083 31708 17132 31736
rect 17083 31705 17095 31708
rect 17037 31699 17095 31705
rect 17126 31696 17132 31708
rect 17184 31696 17190 31748
rect 20162 31736 20168 31748
rect 18262 31708 20168 31736
rect 18800 31680 18828 31708
rect 20162 31696 20168 31708
rect 20220 31696 20226 31748
rect 15933 31671 15991 31677
rect 15933 31637 15945 31671
rect 15979 31668 15991 31671
rect 16666 31668 16672 31680
rect 15979 31640 16672 31668
rect 15979 31637 15991 31640
rect 15933 31631 15991 31637
rect 16666 31628 16672 31640
rect 16724 31628 16730 31680
rect 18782 31628 18788 31680
rect 18840 31628 18846 31680
rect 21634 31628 21640 31680
rect 21692 31628 21698 31680
rect 22002 31628 22008 31680
rect 22060 31628 22066 31680
rect 22370 31628 22376 31680
rect 22428 31668 22434 31680
rect 22646 31668 22652 31680
rect 22428 31640 22652 31668
rect 22428 31628 22434 31640
rect 22646 31628 22652 31640
rect 22704 31668 22710 31680
rect 23385 31671 23443 31677
rect 23385 31668 23397 31671
rect 22704 31640 23397 31668
rect 22704 31628 22710 31640
rect 23385 31637 23397 31640
rect 23431 31637 23443 31671
rect 23385 31631 23443 31637
rect 24026 31628 24032 31680
rect 24084 31628 24090 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 15565 31467 15623 31473
rect 15565 31464 15577 31467
rect 14936 31436 15577 31464
rect 14458 31356 14464 31408
rect 14516 31356 14522 31408
rect 14936 31405 14964 31436
rect 15565 31433 15577 31436
rect 15611 31464 15623 31467
rect 16206 31464 16212 31476
rect 15611 31436 16212 31464
rect 15611 31433 15623 31436
rect 15565 31427 15623 31433
rect 16206 31424 16212 31436
rect 16264 31464 16270 31476
rect 16393 31467 16451 31473
rect 16393 31464 16405 31467
rect 16264 31436 16405 31464
rect 16264 31424 16270 31436
rect 16393 31433 16405 31436
rect 16439 31433 16451 31467
rect 16393 31427 16451 31433
rect 17126 31424 17132 31476
rect 17184 31464 17190 31476
rect 19153 31467 19211 31473
rect 17184 31436 19012 31464
rect 17184 31424 17190 31436
rect 14921 31399 14979 31405
rect 14921 31365 14933 31399
rect 14967 31365 14979 31399
rect 14921 31359 14979 31365
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 17405 31331 17463 31337
rect 17405 31328 17417 31331
rect 16816 31300 17417 31328
rect 16816 31288 16822 31300
rect 17405 31297 17417 31300
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 18782 31288 18788 31340
rect 18840 31288 18846 31340
rect 13538 31220 13544 31272
rect 13596 31260 13602 31272
rect 15197 31263 15255 31269
rect 15197 31260 15209 31263
rect 13596 31232 15209 31260
rect 13596 31220 13602 31232
rect 15197 31229 15209 31232
rect 15243 31260 15255 31263
rect 15470 31260 15476 31272
rect 15243 31232 15476 31260
rect 15243 31229 15255 31232
rect 15197 31223 15255 31229
rect 15470 31220 15476 31232
rect 15528 31220 15534 31272
rect 17681 31263 17739 31269
rect 17681 31229 17693 31263
rect 17727 31260 17739 31263
rect 17770 31260 17776 31272
rect 17727 31232 17776 31260
rect 17727 31229 17739 31232
rect 17681 31223 17739 31229
rect 17770 31220 17776 31232
rect 17828 31220 17834 31272
rect 18984 31260 19012 31436
rect 19153 31433 19165 31467
rect 19199 31464 19211 31467
rect 19702 31464 19708 31476
rect 19199 31436 19708 31464
rect 19199 31433 19211 31436
rect 19153 31427 19211 31433
rect 19702 31424 19708 31436
rect 19760 31424 19766 31476
rect 20533 31467 20591 31473
rect 20533 31433 20545 31467
rect 20579 31464 20591 31467
rect 25498 31464 25504 31476
rect 20579 31436 25504 31464
rect 20579 31433 20591 31436
rect 20533 31427 20591 31433
rect 25498 31424 25504 31436
rect 25556 31424 25562 31476
rect 20162 31356 20168 31408
rect 20220 31396 20226 31408
rect 21269 31399 21327 31405
rect 21269 31396 21281 31399
rect 20220 31368 21281 31396
rect 20220 31356 20226 31368
rect 21269 31365 21281 31368
rect 21315 31365 21327 31399
rect 21269 31359 21327 31365
rect 21545 31399 21603 31405
rect 21545 31365 21557 31399
rect 21591 31396 21603 31399
rect 21726 31396 21732 31408
rect 21591 31368 21732 31396
rect 21591 31365 21603 31368
rect 21545 31359 21603 31365
rect 21726 31356 21732 31368
rect 21784 31396 21790 31408
rect 22002 31396 22008 31408
rect 21784 31368 22008 31396
rect 21784 31356 21790 31368
rect 22002 31356 22008 31368
rect 22060 31396 22066 31408
rect 22060 31356 22094 31396
rect 22646 31356 22652 31408
rect 22704 31396 22710 31408
rect 22741 31399 22799 31405
rect 22741 31396 22753 31399
rect 22704 31368 22753 31396
rect 22704 31356 22710 31368
rect 22741 31365 22753 31368
rect 22787 31396 22799 31399
rect 23014 31396 23020 31408
rect 22787 31368 23020 31396
rect 22787 31365 22799 31368
rect 22741 31359 22799 31365
rect 23014 31356 23020 31368
rect 23072 31356 23078 31408
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31328 19855 31331
rect 20254 31328 20260 31340
rect 19843 31300 20260 31328
rect 19843 31297 19855 31300
rect 19797 31291 19855 31297
rect 20254 31288 20260 31300
rect 20312 31328 20318 31340
rect 20441 31331 20499 31337
rect 20441 31328 20453 31331
rect 20312 31300 20453 31328
rect 20312 31288 20318 31300
rect 20441 31297 20453 31300
rect 20487 31328 20499 31331
rect 21450 31328 21456 31340
rect 20487 31300 21456 31328
rect 20487 31297 20499 31300
rect 20441 31291 20499 31297
rect 21450 31288 21456 31300
rect 21508 31288 21514 31340
rect 20625 31263 20683 31269
rect 20625 31260 20637 31263
rect 18984 31232 20637 31260
rect 20625 31229 20637 31232
rect 20671 31229 20683 31263
rect 20625 31223 20683 31229
rect 20073 31195 20131 31201
rect 20073 31192 20085 31195
rect 18708 31164 20085 31192
rect 13446 31084 13452 31136
rect 13504 31084 13510 31136
rect 14458 31084 14464 31136
rect 14516 31124 14522 31136
rect 15749 31127 15807 31133
rect 15749 31124 15761 31127
rect 14516 31096 15761 31124
rect 14516 31084 14522 31096
rect 15749 31093 15761 31096
rect 15795 31124 15807 31127
rect 16574 31124 16580 31136
rect 15795 31096 16580 31124
rect 15795 31093 15807 31096
rect 15749 31087 15807 31093
rect 16574 31084 16580 31096
rect 16632 31084 16638 31136
rect 16761 31127 16819 31133
rect 16761 31093 16773 31127
rect 16807 31124 16819 31127
rect 16850 31124 16856 31136
rect 16807 31096 16856 31124
rect 16807 31093 16819 31096
rect 16761 31087 16819 31093
rect 16850 31084 16856 31096
rect 16908 31124 16914 31136
rect 17310 31124 17316 31136
rect 16908 31096 17316 31124
rect 16908 31084 16914 31096
rect 17310 31084 17316 31096
rect 17368 31084 17374 31136
rect 17678 31084 17684 31136
rect 17736 31124 17742 31136
rect 18708 31124 18736 31164
rect 20073 31161 20085 31164
rect 20119 31161 20131 31195
rect 20073 31155 20131 31161
rect 17736 31096 18736 31124
rect 17736 31084 17742 31096
rect 18782 31084 18788 31136
rect 18840 31124 18846 31136
rect 19429 31127 19487 31133
rect 19429 31124 19441 31127
rect 18840 31096 19441 31124
rect 18840 31084 18846 31096
rect 19429 31093 19441 31096
rect 19475 31093 19487 31127
rect 22066 31124 22094 31356
rect 22462 31288 22468 31340
rect 22520 31288 22526 31340
rect 24026 31328 24032 31340
rect 23874 31300 24032 31328
rect 24026 31288 24032 31300
rect 24084 31328 24090 31340
rect 25317 31331 25375 31337
rect 24084 31300 24624 31328
rect 24084 31288 24090 31300
rect 22370 31124 22376 31136
rect 22066 31096 22376 31124
rect 19429 31087 19487 31093
rect 22370 31084 22376 31096
rect 22428 31084 22434 31136
rect 23750 31084 23756 31136
rect 23808 31124 23814 31136
rect 24596 31133 24624 31300
rect 25317 31297 25329 31331
rect 25363 31328 25375 31331
rect 25498 31328 25504 31340
rect 25363 31300 25504 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 24213 31127 24271 31133
rect 24213 31124 24225 31127
rect 23808 31096 24225 31124
rect 23808 31084 23814 31096
rect 24213 31093 24225 31096
rect 24259 31093 24271 31127
rect 24213 31087 24271 31093
rect 24581 31127 24639 31133
rect 24581 31093 24593 31127
rect 24627 31124 24639 31127
rect 24670 31124 24676 31136
rect 24627 31096 24676 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 24670 31084 24676 31096
rect 24728 31084 24734 31136
rect 25130 31084 25136 31136
rect 25188 31084 25194 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 9309 30923 9367 30929
rect 9309 30889 9321 30923
rect 9355 30920 9367 30923
rect 10226 30920 10232 30932
rect 9355 30892 10232 30920
rect 9355 30889 9367 30892
rect 9309 30883 9367 30889
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 15657 30923 15715 30929
rect 15657 30889 15669 30923
rect 15703 30920 15715 30923
rect 15841 30923 15899 30929
rect 15841 30920 15853 30923
rect 15703 30892 15853 30920
rect 15703 30889 15715 30892
rect 15657 30883 15715 30889
rect 15841 30889 15853 30892
rect 15887 30920 15899 30923
rect 16298 30920 16304 30932
rect 15887 30892 16304 30920
rect 15887 30889 15899 30892
rect 15841 30883 15899 30889
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9125 30719 9183 30725
rect 9125 30716 9137 30719
rect 8812 30688 9137 30716
rect 8812 30676 8818 30688
rect 9125 30685 9137 30688
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 15286 30676 15292 30728
rect 15344 30716 15350 30728
rect 15672 30716 15700 30883
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 16761 30923 16819 30929
rect 16761 30889 16773 30923
rect 16807 30920 16819 30923
rect 17126 30920 17132 30932
rect 16807 30892 17132 30920
rect 16807 30889 16819 30892
rect 16761 30883 16819 30889
rect 17126 30880 17132 30892
rect 17184 30880 17190 30932
rect 22465 30923 22523 30929
rect 22465 30889 22477 30923
rect 22511 30920 22523 30923
rect 22646 30920 22652 30932
rect 22511 30892 22652 30920
rect 22511 30889 22523 30892
rect 22465 30883 22523 30889
rect 22646 30880 22652 30892
rect 22704 30880 22710 30932
rect 25498 30880 25504 30932
rect 25556 30880 25562 30932
rect 18509 30787 18567 30793
rect 18509 30753 18521 30787
rect 18555 30784 18567 30787
rect 19426 30784 19432 30796
rect 18555 30756 19432 30784
rect 18555 30753 18567 30756
rect 18509 30747 18567 30753
rect 19426 30744 19432 30756
rect 19484 30784 19490 30796
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 19484 30756 20729 30784
rect 19484 30744 19490 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 20717 30747 20775 30753
rect 22370 30744 22376 30796
rect 22428 30784 22434 30796
rect 22646 30784 22652 30796
rect 22428 30756 22652 30784
rect 22428 30744 22434 30756
rect 22646 30744 22652 30756
rect 22704 30744 22710 30796
rect 15344 30688 15700 30716
rect 15344 30676 15350 30688
rect 14553 30651 14611 30657
rect 14553 30617 14565 30651
rect 14599 30648 14611 30651
rect 14826 30648 14832 30660
rect 14599 30620 14832 30648
rect 14599 30617 14611 30620
rect 14553 30611 14611 30617
rect 14826 30608 14832 30620
rect 14884 30608 14890 30660
rect 18233 30651 18291 30657
rect 17802 30620 17908 30648
rect 17880 30580 17908 30620
rect 18233 30617 18245 30651
rect 18279 30648 18291 30651
rect 18279 30620 18460 30648
rect 18279 30617 18291 30620
rect 18233 30611 18291 30617
rect 18432 30592 18460 30620
rect 20898 30608 20904 30660
rect 20956 30648 20962 30660
rect 20993 30651 21051 30657
rect 20993 30648 21005 30651
rect 20956 30620 21005 30648
rect 20956 30608 20962 30620
rect 20993 30617 21005 30620
rect 21039 30617 21051 30651
rect 22218 30620 22324 30648
rect 20993 30611 21051 30617
rect 18322 30580 18328 30592
rect 17880 30552 18328 30580
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 18414 30540 18420 30592
rect 18472 30540 18478 30592
rect 18782 30540 18788 30592
rect 18840 30540 18846 30592
rect 20254 30540 20260 30592
rect 20312 30540 20318 30592
rect 22296 30580 22324 30620
rect 22370 30608 22376 30660
rect 22428 30648 22434 30660
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 22428 30620 24593 30648
rect 22428 30608 22434 30620
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24581 30611 24639 30617
rect 22833 30583 22891 30589
rect 22833 30580 22845 30583
rect 22296 30552 22845 30580
rect 22833 30549 22845 30552
rect 22879 30580 22891 30583
rect 23201 30583 23259 30589
rect 23201 30580 23213 30583
rect 22879 30552 23213 30580
rect 22879 30549 22891 30552
rect 22833 30543 22891 30549
rect 23201 30549 23213 30552
rect 23247 30580 23259 30583
rect 24670 30580 24676 30592
rect 23247 30552 24676 30580
rect 23247 30549 23259 30552
rect 23201 30543 23259 30549
rect 24670 30540 24676 30552
rect 24728 30540 24734 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 20254 30336 20260 30388
rect 20312 30336 20318 30388
rect 11514 30268 11520 30320
rect 11572 30308 11578 30320
rect 11882 30308 11888 30320
rect 11572 30280 11888 30308
rect 11572 30268 11578 30280
rect 11882 30268 11888 30280
rect 11940 30308 11946 30320
rect 15013 30311 15071 30317
rect 11940 30280 12098 30308
rect 11940 30268 11946 30280
rect 15013 30277 15025 30311
rect 15059 30308 15071 30311
rect 15286 30308 15292 30320
rect 15059 30280 15292 30308
rect 15059 30277 15071 30280
rect 15013 30271 15071 30277
rect 15286 30268 15292 30280
rect 15344 30268 15350 30320
rect 19978 30308 19984 30320
rect 15488 30280 19984 30308
rect 8570 30200 8576 30252
rect 8628 30240 8634 30252
rect 8941 30243 8999 30249
rect 8941 30240 8953 30243
rect 8628 30212 8953 30240
rect 8628 30200 8634 30212
rect 8941 30209 8953 30212
rect 8987 30209 8999 30243
rect 8941 30203 8999 30209
rect 13538 30200 13544 30252
rect 13596 30200 13602 30252
rect 12802 30132 12808 30184
rect 12860 30172 12866 30184
rect 13265 30175 13323 30181
rect 13265 30172 13277 30175
rect 12860 30144 13277 30172
rect 12860 30132 12866 30144
rect 13265 30141 13277 30144
rect 13311 30141 13323 30175
rect 13265 30135 13323 30141
rect 13630 30132 13636 30184
rect 13688 30172 13694 30184
rect 14185 30175 14243 30181
rect 14185 30172 14197 30175
rect 13688 30144 14197 30172
rect 13688 30132 13694 30144
rect 14185 30141 14197 30144
rect 14231 30141 14243 30175
rect 14185 30135 14243 30141
rect 14550 30132 14556 30184
rect 14608 30172 14614 30184
rect 15488 30172 15516 30280
rect 19978 30268 19984 30280
rect 20036 30268 20042 30320
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 20530 30308 20536 30320
rect 20395 30280 20536 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 22186 30308 22192 30320
rect 20640 30280 22192 30308
rect 15841 30243 15899 30249
rect 15841 30209 15853 30243
rect 15887 30240 15899 30243
rect 16942 30240 16948 30252
rect 15887 30212 16948 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16942 30200 16948 30212
rect 17000 30200 17006 30252
rect 20640 30240 20668 30280
rect 22186 30268 22192 30280
rect 22244 30268 22250 30320
rect 22465 30311 22523 30317
rect 22465 30277 22477 30311
rect 22511 30308 22523 30311
rect 22738 30308 22744 30320
rect 22511 30280 22744 30308
rect 22511 30277 22523 30280
rect 22465 30271 22523 30277
rect 22738 30268 22744 30280
rect 22796 30268 22802 30320
rect 17052 30212 20668 30240
rect 21453 30243 21511 30249
rect 14608 30144 15516 30172
rect 14608 30132 14614 30144
rect 15562 30132 15568 30184
rect 15620 30132 15626 30184
rect 15749 30175 15807 30181
rect 15749 30141 15761 30175
rect 15795 30172 15807 30175
rect 16758 30172 16764 30184
rect 15795 30144 16764 30172
rect 15795 30141 15807 30144
rect 15749 30135 15807 30141
rect 16758 30132 16764 30144
rect 16816 30172 16822 30184
rect 17052 30172 17080 30212
rect 21453 30209 21465 30243
rect 21499 30240 21511 30243
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21499 30212 22385 30240
rect 21499 30209 21511 30212
rect 21453 30203 21511 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 24670 30200 24676 30252
rect 24728 30200 24734 30252
rect 16816 30144 17080 30172
rect 16816 30132 16822 30144
rect 20438 30132 20444 30184
rect 20496 30132 20502 30184
rect 22554 30132 22560 30184
rect 22612 30132 22618 30184
rect 23290 30132 23296 30184
rect 23348 30132 23354 30184
rect 23569 30175 23627 30181
rect 23569 30141 23581 30175
rect 23615 30172 23627 30175
rect 23658 30172 23664 30184
rect 23615 30144 23664 30172
rect 23615 30141 23627 30144
rect 23569 30135 23627 30141
rect 23658 30132 23664 30144
rect 23716 30132 23722 30184
rect 24854 30132 24860 30184
rect 24912 30172 24918 30184
rect 25041 30175 25099 30181
rect 25041 30172 25053 30175
rect 24912 30144 25053 30172
rect 24912 30132 24918 30144
rect 25041 30141 25053 30144
rect 25087 30141 25099 30175
rect 25041 30135 25099 30141
rect 9030 30064 9036 30116
rect 9088 30104 9094 30116
rect 9125 30107 9183 30113
rect 9125 30104 9137 30107
rect 9088 30076 9137 30104
rect 9088 30064 9094 30076
rect 9125 30073 9137 30076
rect 9171 30073 9183 30107
rect 9125 30067 9183 30073
rect 16298 30064 16304 30116
rect 16356 30104 16362 30116
rect 16356 30076 23428 30104
rect 16356 30064 16362 30076
rect 11790 29996 11796 30048
rect 11848 29996 11854 30048
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 16209 30039 16267 30045
rect 16209 30036 16221 30039
rect 15988 30008 16221 30036
rect 15988 29996 15994 30008
rect 16209 30005 16221 30008
rect 16255 30005 16267 30039
rect 16209 29999 16267 30005
rect 16942 29996 16948 30048
rect 17000 29996 17006 30048
rect 18322 29996 18328 30048
rect 18380 30036 18386 30048
rect 18782 30036 18788 30048
rect 18380 30008 18788 30036
rect 18380 29996 18386 30008
rect 18782 29996 18788 30008
rect 18840 30036 18846 30048
rect 18877 30039 18935 30045
rect 18877 30036 18889 30039
rect 18840 30008 18889 30036
rect 18840 29996 18846 30008
rect 18877 30005 18889 30008
rect 18923 30005 18935 30039
rect 18877 29999 18935 30005
rect 19889 30039 19947 30045
rect 19889 30005 19901 30039
rect 19935 30036 19947 30039
rect 20070 30036 20076 30048
rect 19935 30008 20076 30036
rect 19935 30005 19947 30008
rect 19889 29999 19947 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 21726 29996 21732 30048
rect 21784 30036 21790 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21784 30008 22017 30036
rect 21784 29996 21790 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 23400 30036 23428 30076
rect 26510 30036 26516 30048
rect 23400 30008 26516 30036
rect 22005 29999 22063 30005
rect 26510 29996 26516 30008
rect 26568 29996 26574 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 12802 29792 12808 29844
rect 12860 29832 12866 29844
rect 12897 29835 12955 29841
rect 12897 29832 12909 29835
rect 12860 29804 12909 29832
rect 12860 29792 12866 29804
rect 12897 29801 12909 29804
rect 12943 29801 12955 29835
rect 12897 29795 12955 29801
rect 12912 29764 12940 29795
rect 12986 29792 12992 29844
rect 13044 29832 13050 29844
rect 13446 29832 13452 29844
rect 13044 29804 13452 29832
rect 13044 29792 13050 29804
rect 13446 29792 13452 29804
rect 13504 29792 13510 29844
rect 16298 29792 16304 29844
rect 16356 29792 16362 29844
rect 16942 29792 16948 29844
rect 17000 29832 17006 29844
rect 22094 29832 22100 29844
rect 17000 29804 22100 29832
rect 17000 29792 17006 29804
rect 22094 29792 22100 29804
rect 22152 29792 22158 29844
rect 24578 29792 24584 29844
rect 24636 29792 24642 29844
rect 15562 29764 15568 29776
rect 12912 29736 15568 29764
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11422 29696 11428 29708
rect 11195 29668 11428 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11422 29656 11428 29668
rect 11480 29696 11486 29708
rect 13630 29696 13636 29708
rect 11480 29668 13636 29696
rect 11480 29656 11486 29668
rect 13630 29656 13636 29668
rect 13688 29656 13694 29708
rect 15304 29705 15332 29736
rect 15562 29724 15568 29736
rect 15620 29724 15626 29776
rect 18966 29724 18972 29776
rect 19024 29764 19030 29776
rect 20165 29767 20223 29773
rect 20165 29764 20177 29767
rect 19024 29736 20177 29764
rect 19024 29724 19030 29736
rect 20165 29733 20177 29736
rect 20211 29733 20223 29767
rect 20165 29727 20223 29733
rect 23382 29724 23388 29776
rect 23440 29764 23446 29776
rect 25133 29767 25191 29773
rect 25133 29764 25145 29767
rect 23440 29736 25145 29764
rect 23440 29724 23446 29736
rect 25133 29733 25145 29736
rect 25179 29733 25191 29767
rect 25133 29727 25191 29733
rect 15289 29699 15347 29705
rect 15289 29665 15301 29699
rect 15335 29665 15347 29699
rect 15289 29659 15347 29665
rect 15473 29699 15531 29705
rect 15473 29665 15485 29699
rect 15519 29696 15531 29699
rect 15838 29696 15844 29708
rect 15519 29668 15844 29696
rect 15519 29665 15531 29668
rect 15473 29659 15531 29665
rect 15838 29656 15844 29668
rect 15896 29696 15902 29708
rect 16485 29699 16543 29705
rect 16485 29696 16497 29699
rect 15896 29668 16497 29696
rect 15896 29656 15902 29668
rect 16485 29665 16497 29668
rect 16531 29696 16543 29699
rect 19334 29696 19340 29708
rect 16531 29668 19340 29696
rect 16531 29665 16543 29668
rect 16485 29659 16543 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 20346 29656 20352 29708
rect 20404 29696 20410 29708
rect 20625 29699 20683 29705
rect 20625 29696 20637 29699
rect 20404 29668 20637 29696
rect 20404 29656 20410 29668
rect 20625 29665 20637 29668
rect 20671 29665 20683 29699
rect 20625 29659 20683 29665
rect 20717 29699 20775 29705
rect 20717 29665 20729 29699
rect 20763 29665 20775 29699
rect 20717 29659 20775 29665
rect 15194 29588 15200 29640
rect 15252 29628 15258 29640
rect 15565 29631 15623 29637
rect 15565 29628 15577 29631
rect 15252 29600 15577 29628
rect 15252 29588 15258 29600
rect 15565 29597 15577 29600
rect 15611 29628 15623 29631
rect 16298 29628 16304 29640
rect 15611 29600 16304 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 18785 29631 18843 29637
rect 18785 29597 18797 29631
rect 18831 29628 18843 29631
rect 20438 29628 20444 29640
rect 18831 29600 20444 29628
rect 18831 29597 18843 29600
rect 18785 29591 18843 29597
rect 20438 29588 20444 29600
rect 20496 29588 20502 29640
rect 20732 29628 20760 29659
rect 20548 29600 20760 29628
rect 23385 29631 23443 29637
rect 11054 29520 11060 29572
rect 11112 29560 11118 29572
rect 11425 29563 11483 29569
rect 11425 29560 11437 29563
rect 11112 29532 11437 29560
rect 11112 29520 11118 29532
rect 11425 29529 11437 29532
rect 11471 29529 11483 29563
rect 11882 29560 11888 29572
rect 11425 29523 11483 29529
rect 11808 29532 11888 29560
rect 11808 29492 11836 29532
rect 11882 29520 11888 29532
rect 11940 29520 11946 29572
rect 16574 29520 16580 29572
rect 16632 29560 16638 29572
rect 18509 29563 18567 29569
rect 16632 29532 17342 29560
rect 16632 29520 16638 29532
rect 18509 29529 18521 29563
rect 18555 29560 18567 29563
rect 18874 29560 18880 29572
rect 18555 29532 18880 29560
rect 18555 29529 18567 29532
rect 18509 29523 18567 29529
rect 18874 29520 18880 29532
rect 18932 29560 18938 29572
rect 20548 29560 20576 29600
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 24486 29628 24492 29640
rect 23891 29600 24492 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 18932 29532 20576 29560
rect 22925 29563 22983 29569
rect 18932 29520 18938 29532
rect 22925 29529 22937 29563
rect 22971 29560 22983 29563
rect 23400 29560 23428 29591
rect 24486 29588 24492 29600
rect 24544 29588 24550 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 24854 29560 24860 29572
rect 22971 29532 24860 29560
rect 22971 29529 22983 29532
rect 22925 29523 22983 29529
rect 24854 29520 24860 29532
rect 24912 29520 24918 29572
rect 12710 29492 12716 29504
rect 11808 29464 12716 29492
rect 12710 29452 12716 29464
rect 12768 29492 12774 29504
rect 13173 29495 13231 29501
rect 13173 29492 13185 29495
rect 12768 29464 13185 29492
rect 12768 29452 12774 29464
rect 13173 29461 13185 29464
rect 13219 29492 13231 29495
rect 13633 29495 13691 29501
rect 13633 29492 13645 29495
rect 13219 29464 13645 29492
rect 13219 29461 13231 29464
rect 13173 29455 13231 29461
rect 13633 29461 13645 29464
rect 13679 29461 13691 29495
rect 13633 29455 13691 29461
rect 15933 29495 15991 29501
rect 15933 29461 15945 29495
rect 15979 29492 15991 29495
rect 16022 29492 16028 29504
rect 15979 29464 16028 29492
rect 15979 29461 15991 29464
rect 15933 29455 15991 29461
rect 16022 29452 16028 29464
rect 16080 29452 16086 29504
rect 17037 29495 17095 29501
rect 17037 29461 17049 29495
rect 17083 29492 17095 29495
rect 18414 29492 18420 29504
rect 17083 29464 18420 29492
rect 17083 29461 17095 29464
rect 17037 29455 17095 29461
rect 18414 29452 18420 29464
rect 18472 29452 18478 29504
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19208 29464 19441 29492
rect 19208 29452 19214 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20533 29495 20591 29501
rect 20533 29492 20545 29495
rect 20036 29464 20545 29492
rect 20036 29452 20042 29464
rect 20533 29461 20545 29464
rect 20579 29461 20591 29495
rect 20533 29455 20591 29461
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 23201 29495 23259 29501
rect 23201 29492 23213 29495
rect 22520 29464 23213 29492
rect 22520 29452 22526 29464
rect 23201 29461 23213 29464
rect 23247 29461 23259 29495
rect 23201 29455 23259 29461
rect 24026 29452 24032 29504
rect 24084 29452 24090 29504
rect 24486 29452 24492 29504
rect 24544 29452 24550 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 8846 29248 8852 29300
rect 8904 29288 8910 29300
rect 9493 29291 9551 29297
rect 9493 29288 9505 29291
rect 8904 29260 9505 29288
rect 8904 29248 8910 29260
rect 9493 29257 9505 29260
rect 9539 29257 9551 29291
rect 9493 29251 9551 29257
rect 12526 29248 12532 29300
rect 12584 29248 12590 29300
rect 12618 29248 12624 29300
rect 12676 29248 12682 29300
rect 13538 29248 13544 29300
rect 13596 29288 13602 29300
rect 13596 29260 14044 29288
rect 13596 29248 13602 29260
rect 9953 29223 10011 29229
rect 9953 29189 9965 29223
rect 9999 29220 10011 29223
rect 10226 29220 10232 29232
rect 9999 29192 10232 29220
rect 9999 29189 10011 29192
rect 9953 29183 10011 29189
rect 10226 29180 10232 29192
rect 10284 29180 10290 29232
rect 13630 29220 13636 29232
rect 13372 29192 13636 29220
rect 9861 29155 9919 29161
rect 9861 29121 9873 29155
rect 9907 29152 9919 29155
rect 10410 29152 10416 29164
rect 9907 29124 10416 29152
rect 9907 29121 9919 29124
rect 9861 29115 9919 29121
rect 10410 29112 10416 29124
rect 10468 29112 10474 29164
rect 13372 29161 13400 29192
rect 13630 29180 13636 29192
rect 13688 29180 13694 29232
rect 14016 29220 14044 29260
rect 15102 29248 15108 29300
rect 15160 29248 15166 29300
rect 15930 29248 15936 29300
rect 15988 29248 15994 29300
rect 16022 29248 16028 29300
rect 16080 29248 16086 29300
rect 17313 29291 17371 29297
rect 17313 29257 17325 29291
rect 17359 29288 17371 29291
rect 17402 29288 17408 29300
rect 17359 29260 17408 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 17402 29248 17408 29260
rect 17460 29288 17466 29300
rect 17865 29291 17923 29297
rect 17865 29288 17877 29291
rect 17460 29260 17877 29288
rect 17460 29248 17466 29260
rect 17865 29257 17877 29260
rect 17911 29257 17923 29291
rect 17865 29251 17923 29257
rect 19150 29248 19156 29300
rect 19208 29248 19214 29300
rect 19242 29248 19248 29300
rect 19300 29248 19306 29300
rect 19334 29248 19340 29300
rect 19392 29288 19398 29300
rect 23566 29288 23572 29300
rect 19392 29260 23572 29288
rect 19392 29248 19398 29260
rect 23566 29248 23572 29260
rect 23624 29248 23630 29300
rect 23937 29291 23995 29297
rect 23937 29257 23949 29291
rect 23983 29288 23995 29291
rect 24578 29288 24584 29300
rect 23983 29260 24584 29288
rect 23983 29257 23995 29260
rect 23937 29251 23995 29257
rect 15120 29220 15148 29248
rect 14016 29192 14122 29220
rect 15120 29192 17448 29220
rect 13357 29155 13415 29161
rect 13357 29121 13369 29155
rect 13403 29121 13415 29155
rect 13357 29115 13415 29121
rect 17218 29112 17224 29164
rect 17276 29112 17282 29164
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10045 29087 10103 29093
rect 10045 29084 10057 29087
rect 9732 29056 10057 29084
rect 9732 29044 9738 29056
rect 10045 29053 10057 29056
rect 10091 29053 10103 29087
rect 10045 29047 10103 29053
rect 11514 29044 11520 29096
rect 11572 29084 11578 29096
rect 12805 29087 12863 29093
rect 12805 29084 12817 29087
rect 11572 29056 12817 29084
rect 11572 29044 11578 29056
rect 12805 29053 12817 29056
rect 12851 29084 12863 29087
rect 12986 29084 12992 29096
rect 12851 29056 12992 29084
rect 12851 29053 12863 29056
rect 12805 29047 12863 29053
rect 12986 29044 12992 29056
rect 13044 29044 13050 29096
rect 16117 29087 16175 29093
rect 16117 29084 16129 29087
rect 13464 29056 16129 29084
rect 11974 28976 11980 29028
rect 12032 29016 12038 29028
rect 12161 29019 12219 29025
rect 12161 29016 12173 29019
rect 12032 28988 12173 29016
rect 12032 28976 12038 28988
rect 12161 28985 12173 28988
rect 12207 28985 12219 29019
rect 13464 29016 13492 29056
rect 16117 29053 16129 29056
rect 16163 29053 16175 29087
rect 16117 29047 16175 29053
rect 12161 28979 12219 28985
rect 12406 28988 13492 29016
rect 11330 28908 11336 28960
rect 11388 28948 11394 28960
rect 11790 28948 11796 28960
rect 11388 28920 11796 28948
rect 11388 28908 11394 28920
rect 11790 28908 11796 28920
rect 11848 28948 11854 28960
rect 12406 28948 12434 28988
rect 14642 28976 14648 29028
rect 14700 29016 14706 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 14700 28988 15577 29016
rect 14700 28976 14706 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 15565 28979 15623 28985
rect 15746 28976 15752 29028
rect 15804 29016 15810 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 15804 28988 16865 29016
rect 15804 28976 15810 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 17236 29016 17264 29112
rect 17420 29096 17448 29192
rect 19978 29180 19984 29232
rect 20036 29180 20042 29232
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 19058 29044 19064 29096
rect 19116 29084 19122 29096
rect 19337 29087 19395 29093
rect 19337 29084 19349 29087
rect 19116 29056 19349 29084
rect 19116 29044 19122 29056
rect 19337 29053 19349 29056
rect 19383 29053 19395 29087
rect 19996 29084 20024 29180
rect 21266 29112 21272 29164
rect 21324 29152 21330 29164
rect 21818 29152 21824 29164
rect 21324 29124 21824 29152
rect 21324 29112 21330 29124
rect 21818 29112 21824 29124
rect 21876 29152 21882 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 21876 29124 22201 29152
rect 21876 29112 21882 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 23952 29152 23980 29251
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25409 29291 25467 29297
rect 25409 29288 25421 29291
rect 25372 29260 25421 29288
rect 25372 29248 25378 29260
rect 25409 29257 25421 29260
rect 25455 29257 25467 29291
rect 25409 29251 25467 29257
rect 24946 29180 24952 29232
rect 25004 29220 25010 29232
rect 25498 29220 25504 29232
rect 25004 29192 25504 29220
rect 25004 29180 25010 29192
rect 25498 29180 25504 29192
rect 25556 29180 25562 29232
rect 22189 29115 22247 29121
rect 22940 29124 23980 29152
rect 24029 29155 24087 29161
rect 22940 29084 22968 29124
rect 24029 29121 24041 29155
rect 24075 29152 24087 29155
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 24075 29124 25329 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 25317 29121 25329 29124
rect 25363 29152 25375 29155
rect 26418 29152 26424 29164
rect 25363 29124 26424 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 26418 29112 26424 29124
rect 26476 29112 26482 29164
rect 19996 29056 22968 29084
rect 23017 29087 23075 29093
rect 19337 29047 19395 29053
rect 23017 29053 23029 29087
rect 23063 29084 23075 29087
rect 23290 29084 23296 29096
rect 23063 29056 23296 29084
rect 23063 29053 23075 29056
rect 23017 29047 23075 29053
rect 23290 29044 23296 29056
rect 23348 29084 23354 29096
rect 23474 29084 23480 29096
rect 23348 29056 23480 29084
rect 23348 29044 23354 29056
rect 23474 29044 23480 29056
rect 23532 29044 23538 29096
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 24121 29087 24179 29093
rect 24121 29084 24133 29087
rect 23808 29056 24133 29084
rect 23808 29044 23814 29056
rect 24121 29053 24133 29056
rect 24167 29053 24179 29087
rect 24121 29047 24179 29053
rect 24946 29044 24952 29096
rect 25004 29044 25010 29096
rect 17678 29016 17684 29028
rect 17236 28988 17684 29016
rect 16853 28979 16911 28985
rect 17678 28976 17684 28988
rect 17736 29016 17742 29028
rect 18049 29019 18107 29025
rect 18049 29016 18061 29019
rect 17736 28988 18061 29016
rect 17736 28976 17742 28988
rect 18049 28985 18061 28988
rect 18095 28985 18107 29019
rect 18049 28979 18107 28985
rect 18782 28976 18788 29028
rect 18840 28976 18846 29028
rect 23569 29019 23627 29025
rect 23569 28985 23581 29019
rect 23615 29016 23627 29019
rect 24210 29016 24216 29028
rect 23615 28988 24216 29016
rect 23615 28985 23627 28988
rect 23569 28979 23627 28985
rect 24210 28976 24216 28988
rect 24268 28976 24274 29028
rect 25866 28976 25872 29028
rect 25924 29016 25930 29028
rect 26418 29016 26424 29028
rect 25924 28988 26424 29016
rect 25924 28976 25930 28988
rect 26418 28976 26424 28988
rect 26476 28976 26482 29028
rect 11848 28920 12434 28948
rect 11848 28908 11854 28920
rect 13354 28908 13360 28960
rect 13412 28948 13418 28960
rect 13614 28951 13672 28957
rect 13614 28948 13626 28951
rect 13412 28920 13626 28948
rect 13412 28908 13418 28920
rect 13614 28917 13626 28920
rect 13660 28917 13672 28951
rect 13614 28911 13672 28917
rect 16482 28908 16488 28960
rect 16540 28948 16546 28960
rect 26878 28948 26884 28960
rect 16540 28920 26884 28948
rect 16540 28908 16546 28920
rect 26878 28908 26884 28920
rect 26936 28908 26942 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 9125 28747 9183 28753
rect 9125 28713 9137 28747
rect 9171 28744 9183 28747
rect 9582 28744 9588 28756
rect 9171 28716 9588 28744
rect 9171 28713 9183 28716
rect 9125 28707 9183 28713
rect 9582 28704 9588 28716
rect 9640 28704 9646 28756
rect 18874 28704 18880 28756
rect 18932 28704 18938 28756
rect 22373 28747 22431 28753
rect 22373 28713 22385 28747
rect 22419 28744 22431 28747
rect 23750 28744 23756 28756
rect 22419 28716 23756 28744
rect 22419 28713 22431 28716
rect 22373 28707 22431 28713
rect 23750 28704 23756 28716
rect 23808 28704 23814 28756
rect 21910 28636 21916 28688
rect 21968 28676 21974 28688
rect 22833 28679 22891 28685
rect 22833 28676 22845 28679
rect 21968 28648 22845 28676
rect 21968 28636 21974 28648
rect 22833 28645 22845 28648
rect 22879 28645 22891 28679
rect 22833 28639 22891 28645
rect 22922 28636 22928 28688
rect 22980 28676 22986 28688
rect 25866 28676 25872 28688
rect 22980 28648 25872 28676
rect 22980 28636 22986 28648
rect 25866 28636 25872 28648
rect 25924 28636 25930 28688
rect 15378 28568 15384 28620
rect 15436 28568 15442 28620
rect 15470 28568 15476 28620
rect 15528 28608 15534 28620
rect 15841 28611 15899 28617
rect 15841 28608 15853 28611
rect 15528 28580 15853 28608
rect 15528 28568 15534 28580
rect 15841 28577 15853 28580
rect 15887 28608 15899 28611
rect 16390 28608 16396 28620
rect 15887 28580 16396 28608
rect 15887 28577 15899 28580
rect 15841 28571 15899 28577
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28608 17463 28611
rect 18690 28608 18696 28620
rect 17451 28580 18696 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 18690 28568 18696 28580
rect 18748 28568 18754 28620
rect 20073 28611 20131 28617
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 20898 28608 20904 28620
rect 20119 28580 20904 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 20898 28568 20904 28580
rect 20956 28568 20962 28620
rect 21358 28568 21364 28620
rect 21416 28608 21422 28620
rect 21416 28580 21956 28608
rect 21416 28568 21422 28580
rect 10873 28543 10931 28549
rect 10873 28509 10885 28543
rect 10919 28540 10931 28543
rect 11422 28540 11428 28552
rect 10919 28512 11428 28540
rect 10919 28509 10931 28512
rect 10873 28503 10931 28509
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 14826 28500 14832 28552
rect 14884 28540 14890 28552
rect 17129 28543 17187 28549
rect 17129 28540 17141 28543
rect 14884 28512 17141 28540
rect 14884 28500 14890 28512
rect 17129 28509 17141 28512
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 20438 28500 20444 28552
rect 20496 28540 20502 28552
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 20496 28512 20637 28540
rect 20496 28500 20502 28512
rect 20625 28509 20637 28512
rect 20671 28509 20683 28543
rect 21928 28540 21956 28580
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 23385 28611 23443 28617
rect 23385 28608 23397 28611
rect 22152 28580 23397 28608
rect 22152 28568 22158 28580
rect 23385 28577 23397 28580
rect 23431 28577 23443 28611
rect 23385 28571 23443 28577
rect 25133 28611 25191 28617
rect 25133 28577 25145 28611
rect 25179 28608 25191 28611
rect 25406 28608 25412 28620
rect 25179 28580 25412 28608
rect 25179 28577 25191 28580
rect 25133 28571 25191 28577
rect 25406 28568 25412 28580
rect 25464 28568 25470 28620
rect 23934 28540 23940 28552
rect 21928 28512 23940 28540
rect 20625 28503 20683 28509
rect 23934 28500 23940 28512
rect 23992 28500 23998 28552
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 25041 28543 25099 28549
rect 25041 28509 25053 28543
rect 25087 28540 25099 28543
rect 25222 28540 25228 28552
rect 25087 28512 25228 28540
rect 25087 28509 25099 28512
rect 25041 28503 25099 28509
rect 25222 28500 25228 28512
rect 25280 28500 25286 28552
rect 9582 28432 9588 28484
rect 9640 28432 9646 28484
rect 10597 28475 10655 28481
rect 10597 28441 10609 28475
rect 10643 28472 10655 28475
rect 10962 28472 10968 28484
rect 10643 28444 10968 28472
rect 10643 28441 10655 28444
rect 10597 28435 10655 28441
rect 10962 28432 10968 28444
rect 11020 28432 11026 28484
rect 11330 28432 11336 28484
rect 11388 28472 11394 28484
rect 11701 28475 11759 28481
rect 11701 28472 11713 28475
rect 11388 28444 11713 28472
rect 11388 28432 11394 28444
rect 11701 28441 11713 28444
rect 11747 28441 11759 28475
rect 11701 28435 11759 28441
rect 12710 28432 12716 28484
rect 12768 28432 12774 28484
rect 15289 28475 15347 28481
rect 15289 28441 15301 28475
rect 15335 28472 15347 28475
rect 15335 28444 16344 28472
rect 15335 28441 15347 28444
rect 15289 28435 15347 28441
rect 16316 28416 16344 28444
rect 16390 28432 16396 28484
rect 16448 28472 16454 28484
rect 16448 28444 17894 28472
rect 16448 28432 16454 28444
rect 13173 28407 13231 28413
rect 13173 28373 13185 28407
rect 13219 28404 13231 28407
rect 13354 28404 13360 28416
rect 13219 28376 13360 28404
rect 13219 28373 13231 28376
rect 13173 28367 13231 28373
rect 13354 28364 13360 28376
rect 13412 28364 13418 28416
rect 13538 28364 13544 28416
rect 13596 28364 13602 28416
rect 13814 28364 13820 28416
rect 13872 28404 13878 28416
rect 14829 28407 14887 28413
rect 14829 28404 14841 28407
rect 13872 28376 14841 28404
rect 13872 28364 13878 28376
rect 14829 28373 14841 28376
rect 14875 28373 14887 28407
rect 14829 28367 14887 28373
rect 15197 28407 15255 28413
rect 15197 28373 15209 28407
rect 15243 28404 15255 28407
rect 15562 28404 15568 28416
rect 15243 28376 15568 28404
rect 15243 28373 15255 28376
rect 15197 28367 15255 28373
rect 15562 28364 15568 28376
rect 15620 28364 15626 28416
rect 16114 28364 16120 28416
rect 16172 28364 16178 28416
rect 16298 28364 16304 28416
rect 16356 28364 16362 28416
rect 17788 28404 17816 28444
rect 19058 28432 19064 28484
rect 19116 28472 19122 28484
rect 20901 28475 20959 28481
rect 20901 28472 20913 28475
rect 19116 28444 20913 28472
rect 19116 28432 19122 28444
rect 20901 28441 20913 28444
rect 20947 28441 20959 28475
rect 20901 28435 20959 28441
rect 21358 28432 21364 28484
rect 21416 28432 21422 28484
rect 23293 28475 23351 28481
rect 23293 28441 23305 28475
rect 23339 28472 23351 28475
rect 26050 28472 26056 28484
rect 23339 28444 26056 28472
rect 23339 28441 23351 28444
rect 23293 28435 23351 28441
rect 26050 28432 26056 28444
rect 26108 28432 26114 28484
rect 18322 28404 18328 28416
rect 17788 28376 18328 28404
rect 18322 28364 18328 28376
rect 18380 28364 18386 28416
rect 19429 28407 19487 28413
rect 19429 28373 19441 28407
rect 19475 28404 19487 28407
rect 19518 28404 19524 28416
rect 19475 28376 19524 28404
rect 19475 28373 19487 28376
rect 19429 28367 19487 28373
rect 19518 28364 19524 28376
rect 19576 28364 19582 28416
rect 19794 28364 19800 28416
rect 19852 28364 19858 28416
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 21634 28404 21640 28416
rect 19935 28376 21640 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 22186 28364 22192 28416
rect 22244 28404 22250 28416
rect 22646 28404 22652 28416
rect 22244 28376 22652 28404
rect 22244 28364 22250 28376
rect 22646 28364 22652 28376
rect 22704 28404 22710 28416
rect 23201 28407 23259 28413
rect 23201 28404 23213 28407
rect 22704 28376 23213 28404
rect 22704 28364 22710 28376
rect 23201 28373 23213 28376
rect 23247 28373 23259 28407
rect 23201 28367 23259 28373
rect 23934 28364 23940 28416
rect 23992 28404 23998 28416
rect 24121 28407 24179 28413
rect 24121 28404 24133 28407
rect 23992 28376 24133 28404
rect 23992 28364 23998 28376
rect 24121 28373 24133 28376
rect 24167 28404 24179 28407
rect 24394 28404 24400 28416
rect 24167 28376 24400 28404
rect 24167 28373 24179 28376
rect 24121 28367 24179 28373
rect 24394 28364 24400 28376
rect 24452 28364 24458 28416
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 24544 28376 24593 28404
rect 24544 28364 24550 28376
rect 24581 28373 24593 28376
rect 24627 28373 24639 28407
rect 24581 28367 24639 28373
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 12710 28200 12716 28212
rect 12406 28172 12716 28200
rect 11057 28135 11115 28141
rect 11057 28101 11069 28135
rect 11103 28132 11115 28135
rect 12406 28132 12434 28172
rect 12710 28160 12716 28172
rect 12768 28200 12774 28212
rect 13538 28200 13544 28212
rect 12768 28172 13544 28200
rect 12768 28160 12774 28172
rect 13538 28160 13544 28172
rect 13596 28200 13602 28212
rect 13725 28203 13783 28209
rect 13725 28200 13737 28203
rect 13596 28172 13737 28200
rect 13596 28160 13602 28172
rect 13725 28169 13737 28172
rect 13771 28169 13783 28203
rect 13725 28163 13783 28169
rect 15565 28203 15623 28209
rect 15565 28169 15577 28203
rect 15611 28200 15623 28203
rect 16390 28200 16396 28212
rect 15611 28172 16396 28200
rect 15611 28169 15623 28172
rect 15565 28163 15623 28169
rect 16390 28160 16396 28172
rect 16448 28200 16454 28212
rect 16485 28203 16543 28209
rect 16485 28200 16497 28203
rect 16448 28172 16497 28200
rect 16448 28160 16454 28172
rect 16485 28169 16497 28172
rect 16531 28200 16543 28203
rect 16531 28172 18736 28200
rect 16531 28169 16543 28172
rect 16485 28163 16543 28169
rect 11103 28104 12466 28132
rect 11103 28101 11115 28104
rect 11057 28095 11115 28101
rect 16666 28092 16672 28144
rect 16724 28132 16730 28144
rect 17221 28135 17279 28141
rect 17221 28132 17233 28135
rect 16724 28104 17233 28132
rect 16724 28092 16730 28104
rect 17221 28101 17233 28104
rect 17267 28132 17279 28135
rect 18598 28132 18604 28144
rect 17267 28104 18604 28132
rect 17267 28101 17279 28104
rect 17221 28095 17279 28101
rect 18598 28092 18604 28104
rect 18656 28092 18662 28144
rect 18708 28132 18736 28172
rect 19794 28160 19800 28212
rect 19852 28200 19858 28212
rect 19889 28203 19947 28209
rect 19889 28200 19901 28203
rect 19852 28172 19901 28200
rect 19852 28160 19858 28172
rect 19889 28169 19901 28172
rect 19935 28169 19947 28203
rect 19889 28163 19947 28169
rect 22465 28203 22523 28209
rect 22465 28169 22477 28203
rect 22511 28200 22523 28203
rect 26234 28200 26240 28212
rect 22511 28172 26240 28200
rect 22511 28169 22523 28172
rect 22465 28163 22523 28169
rect 26234 28160 26240 28172
rect 26292 28160 26298 28212
rect 18708 28104 20668 28132
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28064 15715 28067
rect 16301 28067 16359 28073
rect 16301 28064 16313 28067
rect 15703 28036 16313 28064
rect 15703 28033 15715 28036
rect 15657 28027 15715 28033
rect 16301 28033 16313 28036
rect 16347 28064 16359 28067
rect 16482 28064 16488 28076
rect 16347 28036 16488 28064
rect 16347 28033 16359 28036
rect 16301 28027 16359 28033
rect 16482 28024 16488 28036
rect 16540 28024 16546 28076
rect 17310 28024 17316 28076
rect 17368 28064 17374 28076
rect 18506 28064 18512 28076
rect 17368 28036 18512 28064
rect 17368 28024 17374 28036
rect 18506 28024 18512 28036
rect 18564 28024 18570 28076
rect 11701 27999 11759 28005
rect 11701 27965 11713 27999
rect 11747 27965 11759 27999
rect 11701 27959 11759 27965
rect 11977 27999 12035 28005
rect 11977 27965 11989 27999
rect 12023 27996 12035 27999
rect 12066 27996 12072 28008
rect 12023 27968 12072 27996
rect 12023 27965 12035 27968
rect 11977 27959 12035 27965
rect 9858 27888 9864 27940
rect 9916 27928 9922 27940
rect 11716 27928 11744 27959
rect 12066 27956 12072 27968
rect 12124 27956 12130 28008
rect 13446 27956 13452 28008
rect 13504 27996 13510 28008
rect 15378 27996 15384 28008
rect 13504 27968 15384 27996
rect 13504 27956 13510 27968
rect 15378 27956 15384 27968
rect 15436 27996 15442 28008
rect 15749 27999 15807 28005
rect 15436 27968 15608 27996
rect 15436 27956 15442 27968
rect 14826 27928 14832 27940
rect 9916 27900 11744 27928
rect 9916 27888 9922 27900
rect 11716 27860 11744 27900
rect 13372 27900 14832 27928
rect 13372 27860 13400 27900
rect 14826 27888 14832 27900
rect 14884 27888 14890 27940
rect 15580 27928 15608 27968
rect 15749 27965 15761 27999
rect 15795 27965 15807 27999
rect 15749 27959 15807 27965
rect 15764 27928 15792 27959
rect 17402 27956 17408 28008
rect 17460 27956 17466 28008
rect 17954 27956 17960 28008
rect 18012 27996 18018 28008
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 18012 27968 18061 27996
rect 18012 27956 18018 27968
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 18322 27956 18328 28008
rect 18380 27996 18386 28008
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 18380 27968 18981 27996
rect 18380 27956 18386 27968
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 20438 27956 20444 28008
rect 20496 27956 20502 28008
rect 20640 27996 20668 28104
rect 20806 28092 20812 28144
rect 20864 28132 20870 28144
rect 21358 28132 21364 28144
rect 20864 28104 21364 28132
rect 20864 28092 20870 28104
rect 21358 28092 21364 28104
rect 21416 28092 21422 28144
rect 21542 28092 21548 28144
rect 21600 28132 21606 28144
rect 22373 28135 22431 28141
rect 22373 28132 22385 28135
rect 21600 28104 22385 28132
rect 21600 28092 21606 28104
rect 22373 28101 22385 28104
rect 22419 28132 22431 28135
rect 22554 28132 22560 28144
rect 22419 28104 22560 28132
rect 22419 28101 22431 28104
rect 22373 28095 22431 28101
rect 22554 28092 22560 28104
rect 22612 28132 22618 28144
rect 22922 28132 22928 28144
rect 22612 28104 22928 28132
rect 22612 28092 22618 28104
rect 22922 28092 22928 28104
rect 22980 28092 22986 28144
rect 24394 28132 24400 28144
rect 24242 28104 24400 28132
rect 24394 28092 24400 28104
rect 24452 28132 24458 28144
rect 24670 28132 24676 28144
rect 24452 28104 24676 28132
rect 24452 28092 24458 28104
rect 24670 28092 24676 28104
rect 24728 28132 24734 28144
rect 24946 28132 24952 28144
rect 24728 28104 24952 28132
rect 24728 28092 24734 28104
rect 24946 28092 24952 28104
rect 25004 28132 25010 28144
rect 25225 28135 25283 28141
rect 25225 28132 25237 28135
rect 25004 28104 25237 28132
rect 25004 28092 25010 28104
rect 25225 28101 25237 28104
rect 25271 28101 25283 28135
rect 25225 28095 25283 28101
rect 21266 28024 21272 28076
rect 21324 28024 21330 28076
rect 20640 27968 22094 27996
rect 15580 27900 15792 27928
rect 16666 27888 16672 27940
rect 16724 27928 16730 27940
rect 17034 27928 17040 27940
rect 16724 27900 17040 27928
rect 16724 27888 16730 27900
rect 17034 27888 17040 27900
rect 17092 27928 17098 27940
rect 19337 27931 19395 27937
rect 19337 27928 19349 27931
rect 17092 27900 19349 27928
rect 17092 27888 17098 27900
rect 19337 27897 19349 27900
rect 19383 27928 19395 27931
rect 21266 27928 21272 27940
rect 19383 27900 21272 27928
rect 19383 27897 19395 27900
rect 19337 27891 19395 27897
rect 21266 27888 21272 27900
rect 21324 27888 21330 27940
rect 22066 27928 22094 27968
rect 22554 27956 22560 28008
rect 22612 27956 22618 28008
rect 24118 27996 24124 28008
rect 22664 27968 24124 27996
rect 22664 27928 22692 27968
rect 24118 27956 24124 27968
rect 24176 27956 24182 28008
rect 24670 27956 24676 28008
rect 24728 27956 24734 28008
rect 24949 27999 25007 28005
rect 24949 27965 24961 27999
rect 24995 27965 25007 27999
rect 24949 27959 25007 27965
rect 22066 27900 22692 27928
rect 11716 27832 13400 27860
rect 13446 27820 13452 27872
rect 13504 27820 13510 27872
rect 13906 27820 13912 27872
rect 13964 27860 13970 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 13964 27832 15209 27860
rect 13964 27820 13970 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 16850 27820 16856 27872
rect 16908 27820 16914 27872
rect 18506 27820 18512 27872
rect 18564 27820 18570 27872
rect 18598 27820 18604 27872
rect 18656 27860 18662 27872
rect 18693 27863 18751 27869
rect 18693 27860 18705 27863
rect 18656 27832 18705 27860
rect 18656 27820 18662 27832
rect 18693 27829 18705 27832
rect 18739 27829 18751 27863
rect 18693 27823 18751 27829
rect 21542 27820 21548 27872
rect 21600 27820 21606 27872
rect 21634 27820 21640 27872
rect 21692 27860 21698 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 21692 27832 22017 27860
rect 21692 27820 21698 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 22738 27820 22744 27872
rect 22796 27860 22802 27872
rect 23201 27863 23259 27869
rect 23201 27860 23213 27863
rect 22796 27832 23213 27860
rect 22796 27820 22802 27832
rect 23201 27829 23213 27832
rect 23247 27860 23259 27863
rect 23382 27860 23388 27872
rect 23247 27832 23388 27860
rect 23247 27829 23259 27832
rect 23201 27823 23259 27829
rect 23382 27820 23388 27832
rect 23440 27820 23446 27872
rect 23566 27820 23572 27872
rect 23624 27860 23630 27872
rect 24964 27860 24992 27959
rect 23624 27832 24992 27860
rect 23624 27820 23630 27832
rect 25406 27820 25412 27872
rect 25464 27820 25470 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 11995 27659 12053 27665
rect 11995 27625 12007 27659
rect 12041 27656 12053 27659
rect 13446 27656 13452 27668
rect 12041 27628 13452 27656
rect 12041 27625 12053 27628
rect 11995 27619 12053 27625
rect 13446 27616 13452 27628
rect 13504 27616 13510 27668
rect 21379 27659 21437 27665
rect 21379 27625 21391 27659
rect 21425 27656 21437 27659
rect 22094 27656 22100 27668
rect 21425 27628 22100 27656
rect 21425 27625 21437 27628
rect 21379 27619 21437 27625
rect 22094 27616 22100 27628
rect 22152 27616 22158 27668
rect 23382 27616 23388 27668
rect 23440 27656 23446 27668
rect 23581 27659 23639 27665
rect 23581 27656 23593 27659
rect 23440 27628 23593 27656
rect 23440 27616 23446 27628
rect 23581 27625 23593 27628
rect 23627 27625 23639 27659
rect 23581 27619 23639 27625
rect 12342 27548 12348 27600
rect 12400 27588 12406 27600
rect 12710 27588 12716 27600
rect 12400 27560 12716 27588
rect 12400 27548 12406 27560
rect 12710 27548 12716 27560
rect 12768 27548 12774 27600
rect 24670 27548 24676 27600
rect 24728 27588 24734 27600
rect 24728 27560 25176 27588
rect 24728 27548 24734 27560
rect 11422 27480 11428 27532
rect 11480 27520 11486 27532
rect 12253 27523 12311 27529
rect 12253 27520 12265 27523
rect 11480 27492 12265 27520
rect 11480 27480 11486 27492
rect 12253 27489 12265 27492
rect 12299 27489 12311 27523
rect 13541 27523 13599 27529
rect 13541 27520 13553 27523
rect 12253 27483 12311 27489
rect 12406 27492 13553 27520
rect 11238 27344 11244 27396
rect 11296 27344 11302 27396
rect 9306 27276 9312 27328
rect 9364 27316 9370 27328
rect 10505 27319 10563 27325
rect 10505 27316 10517 27319
rect 9364 27288 10517 27316
rect 9364 27276 9370 27288
rect 10505 27285 10517 27288
rect 10551 27316 10563 27319
rect 12406 27316 12434 27492
rect 13541 27489 13553 27492
rect 13587 27489 13599 27523
rect 13541 27483 13599 27489
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27520 15899 27523
rect 16206 27520 16212 27532
rect 15887 27492 16212 27520
rect 15887 27489 15899 27492
rect 15841 27483 15899 27489
rect 16206 27480 16212 27492
rect 16264 27480 16270 27532
rect 17770 27480 17776 27532
rect 17828 27520 17834 27532
rect 18049 27523 18107 27529
rect 18049 27520 18061 27523
rect 17828 27492 18061 27520
rect 17828 27480 17834 27492
rect 18049 27489 18061 27492
rect 18095 27489 18107 27523
rect 18049 27483 18107 27489
rect 21637 27523 21695 27529
rect 21637 27489 21649 27523
rect 21683 27520 21695 27523
rect 23566 27520 23572 27532
rect 21683 27492 23572 27520
rect 21683 27489 21695 27492
rect 21637 27483 21695 27489
rect 23566 27480 23572 27492
rect 23624 27520 23630 27532
rect 23845 27523 23903 27529
rect 23845 27520 23857 27523
rect 23624 27492 23857 27520
rect 23624 27480 23630 27492
rect 23845 27489 23857 27492
rect 23891 27489 23903 27523
rect 23845 27483 23903 27489
rect 25038 27480 25044 27532
rect 25096 27480 25102 27532
rect 25148 27529 25176 27560
rect 25133 27523 25191 27529
rect 25133 27489 25145 27523
rect 25179 27489 25191 27523
rect 25133 27483 25191 27489
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27452 12679 27455
rect 12710 27452 12716 27464
rect 12667 27424 12716 27452
rect 12667 27421 12679 27424
rect 12621 27415 12679 27421
rect 12710 27412 12716 27424
rect 12768 27412 12774 27464
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 13814 27452 13820 27464
rect 13495 27424 13820 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 14918 27412 14924 27464
rect 14976 27452 14982 27464
rect 16758 27452 16764 27464
rect 14976 27424 16764 27452
rect 14976 27412 14982 27424
rect 16758 27412 16764 27424
rect 16816 27412 16822 27464
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 17954 27452 17960 27464
rect 17911 27424 17960 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 24213 27455 24271 27461
rect 24213 27421 24225 27455
rect 24259 27452 24271 27455
rect 24259 27424 24716 27452
rect 24259 27421 24271 27424
rect 24213 27415 24271 27421
rect 13357 27387 13415 27393
rect 13357 27353 13369 27387
rect 13403 27384 13415 27387
rect 13906 27384 13912 27396
rect 13403 27356 13912 27384
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 13906 27344 13912 27356
rect 13964 27344 13970 27396
rect 15657 27387 15715 27393
rect 15657 27353 15669 27387
rect 15703 27384 15715 27387
rect 15703 27356 16344 27384
rect 15703 27353 15715 27356
rect 15657 27347 15715 27353
rect 16316 27328 16344 27356
rect 20806 27344 20812 27396
rect 20864 27344 20870 27396
rect 22002 27344 22008 27396
rect 22060 27384 22066 27396
rect 24688 27384 24716 27424
rect 24854 27412 24860 27464
rect 24912 27452 24918 27464
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 24912 27424 24961 27452
rect 24912 27412 24918 27424
rect 24949 27421 24961 27424
rect 24995 27452 25007 27455
rect 25406 27452 25412 27464
rect 24995 27424 25412 27452
rect 24995 27421 25007 27424
rect 24949 27415 25007 27421
rect 25406 27412 25412 27424
rect 25464 27412 25470 27464
rect 26050 27384 26056 27396
rect 22060 27356 22402 27384
rect 23216 27356 24624 27384
rect 24688 27356 26056 27384
rect 22060 27344 22066 27356
rect 10551 27288 12434 27316
rect 10551 27285 10563 27288
rect 10505 27279 10563 27285
rect 12618 27276 12624 27328
rect 12676 27316 12682 27328
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12676 27288 13001 27316
rect 12676 27276 12682 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13538 27276 13544 27328
rect 13596 27316 13602 27328
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 13596 27288 15209 27316
rect 13596 27276 13602 27288
rect 15197 27285 15209 27288
rect 15243 27285 15255 27319
rect 15197 27279 15255 27285
rect 15562 27276 15568 27328
rect 15620 27316 15626 27328
rect 16114 27316 16120 27328
rect 15620 27288 16120 27316
rect 15620 27276 15626 27288
rect 16114 27276 16120 27288
rect 16172 27316 16178 27328
rect 16209 27319 16267 27325
rect 16209 27316 16221 27319
rect 16172 27288 16221 27316
rect 16172 27276 16178 27288
rect 16209 27285 16221 27288
rect 16255 27285 16267 27319
rect 16209 27279 16267 27285
rect 16298 27276 16304 27328
rect 16356 27316 16362 27328
rect 16393 27319 16451 27325
rect 16393 27316 16405 27319
rect 16356 27288 16405 27316
rect 16356 27276 16362 27288
rect 16393 27285 16405 27288
rect 16439 27285 16451 27319
rect 16393 27279 16451 27285
rect 16482 27276 16488 27328
rect 16540 27316 16546 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 16540 27288 17509 27316
rect 16540 27276 16546 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 17497 27279 17555 27285
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 17957 27319 18015 27325
rect 17957 27316 17969 27319
rect 17644 27288 17969 27316
rect 17644 27276 17650 27288
rect 17957 27285 17969 27288
rect 18003 27285 18015 27319
rect 17957 27279 18015 27285
rect 19889 27319 19947 27325
rect 19889 27285 19901 27319
rect 19935 27316 19947 27319
rect 20714 27316 20720 27328
rect 19935 27288 20720 27316
rect 19935 27285 19947 27288
rect 19889 27279 19947 27285
rect 20714 27276 20720 27288
rect 20772 27276 20778 27328
rect 22646 27276 22652 27328
rect 22704 27316 22710 27328
rect 23216 27316 23244 27356
rect 24596 27325 24624 27356
rect 26050 27344 26056 27356
rect 26108 27344 26114 27396
rect 22704 27288 23244 27316
rect 24581 27319 24639 27325
rect 22704 27276 22710 27288
rect 24581 27285 24593 27319
rect 24627 27285 24639 27319
rect 24581 27279 24639 27285
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 9582 27072 9588 27124
rect 9640 27112 9646 27124
rect 9640 27084 10916 27112
rect 9640 27072 9646 27084
rect 9858 27044 9864 27056
rect 9324 27016 9864 27044
rect 9324 26985 9352 27016
rect 9858 27004 9864 27016
rect 9916 27004 9922 27056
rect 10888 27044 10916 27084
rect 11054 27072 11060 27124
rect 11112 27072 11118 27124
rect 15657 27115 15715 27121
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16850 27112 16856 27124
rect 15703 27084 16856 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 21542 27112 21548 27124
rect 16960 27084 21548 27112
rect 11238 27044 11244 27056
rect 10810 27016 11244 27044
rect 11238 27004 11244 27016
rect 11296 27004 11302 27056
rect 12710 27004 12716 27056
rect 12768 27044 12774 27056
rect 14553 27047 14611 27053
rect 12768 27016 13386 27044
rect 12768 27004 12774 27016
rect 14553 27013 14565 27047
rect 14599 27044 14611 27047
rect 15102 27044 15108 27056
rect 14599 27016 15108 27044
rect 14599 27013 14611 27016
rect 14553 27007 14611 27013
rect 15102 27004 15108 27016
rect 15160 27004 15166 27056
rect 15746 27004 15752 27056
rect 15804 27004 15810 27056
rect 15930 27004 15936 27056
rect 15988 27044 15994 27056
rect 16960 27044 16988 27084
rect 21542 27072 21548 27084
rect 21600 27072 21606 27124
rect 22370 27072 22376 27124
rect 22428 27112 22434 27124
rect 22741 27115 22799 27121
rect 22741 27112 22753 27115
rect 22428 27084 22753 27112
rect 22428 27072 22434 27084
rect 22741 27081 22753 27084
rect 22787 27081 22799 27115
rect 22741 27075 22799 27081
rect 22830 27072 22836 27124
rect 22888 27072 22894 27124
rect 23658 27112 23664 27124
rect 23032 27084 23664 27112
rect 15988 27016 16988 27044
rect 19429 27047 19487 27053
rect 15988 27004 15994 27016
rect 19429 27013 19441 27047
rect 19475 27044 19487 27047
rect 22094 27044 22100 27056
rect 19475 27016 22100 27044
rect 19475 27013 19487 27016
rect 19429 27007 19487 27013
rect 22094 27004 22100 27016
rect 22152 27044 22158 27056
rect 22554 27044 22560 27056
rect 22152 27016 22560 27044
rect 22152 27004 22158 27016
rect 22554 27004 22560 27016
rect 22612 27004 22618 27056
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26945 9367 26979
rect 9309 26939 9367 26945
rect 14826 26936 14832 26988
rect 14884 26936 14890 26988
rect 18322 26936 18328 26988
rect 18380 26936 18386 26988
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 22370 26976 22376 26988
rect 22244 26948 22376 26976
rect 22244 26936 22250 26948
rect 22370 26936 22376 26948
rect 22428 26936 22434 26988
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 9324 26880 9597 26908
rect 9324 26852 9352 26880
rect 9585 26877 9597 26880
rect 9631 26877 9643 26911
rect 15841 26911 15899 26917
rect 15841 26908 15853 26911
rect 9585 26871 9643 26877
rect 13188 26880 15853 26908
rect 9306 26800 9312 26852
rect 9364 26800 9370 26852
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 11517 26775 11575 26781
rect 11517 26772 11529 26775
rect 11296 26744 11529 26772
rect 11296 26732 11302 26744
rect 11517 26741 11529 26744
rect 11563 26772 11575 26775
rect 12342 26772 12348 26784
rect 11563 26744 12348 26772
rect 11563 26741 11575 26744
rect 11517 26735 11575 26741
rect 12342 26732 12348 26744
rect 12400 26732 12406 26784
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 13081 26775 13139 26781
rect 13081 26772 13093 26775
rect 12584 26744 13093 26772
rect 12584 26732 12590 26744
rect 13081 26741 13093 26744
rect 13127 26772 13139 26775
rect 13188 26772 13216 26880
rect 15841 26877 15853 26880
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 19705 26911 19763 26917
rect 19705 26877 19717 26911
rect 19751 26908 19763 26911
rect 20438 26908 20444 26920
rect 19751 26880 20444 26908
rect 19751 26877 19763 26880
rect 19705 26871 19763 26877
rect 13127 26744 13216 26772
rect 13127 26741 13139 26744
rect 13081 26735 13139 26741
rect 15010 26732 15016 26784
rect 15068 26772 15074 26784
rect 15289 26775 15347 26781
rect 15289 26772 15301 26775
rect 15068 26744 15301 26772
rect 15068 26732 15074 26744
rect 15289 26741 15301 26744
rect 15335 26741 15347 26775
rect 15289 26735 15347 26741
rect 17957 26775 18015 26781
rect 17957 26741 17969 26775
rect 18003 26772 18015 26775
rect 18690 26772 18696 26784
rect 18003 26744 18696 26772
rect 18003 26741 18015 26744
rect 17957 26735 18015 26741
rect 18690 26732 18696 26744
rect 18748 26732 18754 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 19720 26772 19748 26871
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 23032 26917 23060 27084
rect 23658 27072 23664 27084
rect 23716 27072 23722 27124
rect 24670 27072 24676 27124
rect 24728 27112 24734 27124
rect 25317 27115 25375 27121
rect 25317 27112 25329 27115
rect 24728 27084 25329 27112
rect 24728 27072 24734 27084
rect 25317 27081 25329 27084
rect 25363 27081 25375 27115
rect 25317 27075 25375 27081
rect 24946 26936 24952 26988
rect 25004 26936 25010 26988
rect 23017 26911 23075 26917
rect 23017 26877 23029 26911
rect 23063 26877 23075 26911
rect 23017 26871 23075 26877
rect 23566 26868 23572 26920
rect 23624 26868 23630 26920
rect 23845 26911 23903 26917
rect 23845 26877 23857 26911
rect 23891 26908 23903 26911
rect 25406 26908 25412 26920
rect 23891 26880 25412 26908
rect 23891 26877 23903 26880
rect 23845 26871 23903 26877
rect 25406 26868 25412 26880
rect 25464 26868 25470 26920
rect 21266 26800 21272 26852
rect 21324 26840 21330 26852
rect 22373 26843 22431 26849
rect 22373 26840 22385 26843
rect 21324 26812 22385 26840
rect 21324 26800 21330 26812
rect 22373 26809 22385 26812
rect 22419 26809 22431 26843
rect 22373 26803 22431 26809
rect 19484 26744 19748 26772
rect 20073 26775 20131 26781
rect 19484 26732 19490 26744
rect 20073 26741 20085 26775
rect 20119 26772 20131 26775
rect 20162 26772 20168 26784
rect 20119 26744 20168 26772
rect 20119 26741 20131 26744
rect 20073 26735 20131 26741
rect 20162 26732 20168 26744
rect 20220 26772 20226 26784
rect 20806 26772 20812 26784
rect 20220 26744 20812 26772
rect 20220 26732 20226 26744
rect 20806 26732 20812 26744
rect 20864 26772 20870 26784
rect 21821 26775 21879 26781
rect 21821 26772 21833 26775
rect 20864 26744 21833 26772
rect 20864 26732 20870 26744
rect 21821 26741 21833 26744
rect 21867 26772 21879 26775
rect 22002 26772 22008 26784
rect 21867 26744 22008 26772
rect 21867 26741 21879 26744
rect 21821 26735 21879 26741
rect 22002 26732 22008 26744
rect 22060 26732 22066 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 9398 26528 9404 26580
rect 9456 26568 9462 26580
rect 10873 26571 10931 26577
rect 9456 26540 10456 26568
rect 9456 26528 9462 26540
rect 10428 26500 10456 26540
rect 10873 26537 10885 26571
rect 10919 26568 10931 26571
rect 12066 26568 12072 26580
rect 10919 26540 12072 26568
rect 10919 26537 10931 26540
rect 10873 26531 10931 26537
rect 12066 26528 12072 26540
rect 12124 26528 12130 26580
rect 13630 26528 13636 26580
rect 13688 26568 13694 26580
rect 15657 26571 15715 26577
rect 15657 26568 15669 26571
rect 13688 26540 15669 26568
rect 13688 26528 13694 26540
rect 15657 26537 15669 26540
rect 15703 26537 15715 26571
rect 15657 26531 15715 26537
rect 16390 26528 16396 26580
rect 16448 26568 16454 26580
rect 17218 26568 17224 26580
rect 16448 26540 17224 26568
rect 16448 26528 16454 26540
rect 17218 26528 17224 26540
rect 17276 26528 17282 26580
rect 21177 26571 21235 26577
rect 21177 26537 21189 26571
rect 21223 26568 21235 26571
rect 22094 26568 22100 26580
rect 21223 26540 22100 26568
rect 21223 26537 21235 26540
rect 21177 26531 21235 26537
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 24029 26571 24087 26577
rect 24029 26537 24041 26571
rect 24075 26568 24087 26571
rect 24946 26568 24952 26580
rect 24075 26540 24952 26568
rect 24075 26537 24087 26540
rect 24029 26531 24087 26537
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 11333 26503 11391 26509
rect 11333 26500 11345 26503
rect 10428 26472 11345 26500
rect 11333 26469 11345 26472
rect 11379 26500 11391 26503
rect 11514 26500 11520 26512
rect 11379 26472 11520 26500
rect 11379 26469 11391 26472
rect 11333 26463 11391 26469
rect 11514 26460 11520 26472
rect 11572 26460 11578 26512
rect 11606 26460 11612 26512
rect 11664 26500 11670 26512
rect 14277 26503 14335 26509
rect 14277 26500 14289 26503
rect 11664 26472 14289 26500
rect 11664 26460 11670 26472
rect 14277 26469 14289 26472
rect 14323 26469 14335 26503
rect 16574 26500 16580 26512
rect 14277 26463 14335 26469
rect 16132 26472 16580 26500
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 9858 26432 9864 26444
rect 9171 26404 9864 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 9858 26392 9864 26404
rect 9916 26392 9922 26444
rect 14734 26392 14740 26444
rect 14792 26432 14798 26444
rect 14829 26435 14887 26441
rect 14829 26432 14841 26435
rect 14792 26404 14841 26432
rect 14792 26392 14798 26404
rect 14829 26401 14841 26404
rect 14875 26401 14887 26435
rect 14829 26395 14887 26401
rect 15381 26435 15439 26441
rect 15381 26401 15393 26435
rect 15427 26432 15439 26435
rect 15470 26432 15476 26444
rect 15427 26404 15476 26432
rect 15427 26401 15439 26404
rect 15381 26395 15439 26401
rect 15470 26392 15476 26404
rect 15528 26392 15534 26444
rect 16132 26441 16160 26472
rect 16574 26460 16580 26472
rect 16632 26500 16638 26512
rect 17037 26503 17095 26509
rect 17037 26500 17049 26503
rect 16632 26472 17049 26500
rect 16632 26460 16638 26472
rect 17037 26469 17049 26472
rect 17083 26500 17095 26503
rect 17126 26500 17132 26512
rect 17083 26472 17132 26500
rect 17083 26469 17095 26472
rect 17037 26463 17095 26469
rect 17126 26460 17132 26472
rect 17184 26460 17190 26512
rect 20806 26460 20812 26512
rect 20864 26500 20870 26512
rect 21453 26503 21511 26509
rect 21453 26500 21465 26503
rect 20864 26472 21465 26500
rect 20864 26460 20870 26472
rect 21453 26469 21465 26472
rect 21499 26469 21511 26503
rect 21453 26463 21511 26469
rect 22554 26460 22560 26512
rect 22612 26500 22618 26512
rect 22649 26503 22707 26509
rect 22649 26500 22661 26503
rect 22612 26472 22661 26500
rect 22612 26460 22618 26472
rect 22649 26469 22661 26472
rect 22695 26469 22707 26503
rect 22649 26463 22707 26469
rect 24581 26503 24639 26509
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 25222 26500 25228 26512
rect 24627 26472 25228 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 25222 26460 25228 26472
rect 25280 26460 25286 26512
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 16206 26392 16212 26444
rect 16264 26392 16270 26444
rect 16758 26392 16764 26444
rect 16816 26392 16822 26444
rect 16942 26392 16948 26444
rect 17000 26392 17006 26444
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26432 19763 26435
rect 20714 26432 20720 26444
rect 19751 26404 20720 26432
rect 19751 26401 19763 26404
rect 19705 26395 19763 26401
rect 20714 26392 20720 26404
rect 20772 26392 20778 26444
rect 22278 26392 22284 26444
rect 22336 26432 22342 26444
rect 23201 26435 23259 26441
rect 23201 26432 23213 26435
rect 22336 26404 23213 26432
rect 22336 26392 22342 26404
rect 23201 26401 23213 26404
rect 23247 26401 23259 26435
rect 23201 26395 23259 26401
rect 25038 26392 25044 26444
rect 25096 26432 25102 26444
rect 25133 26435 25191 26441
rect 25133 26432 25145 26435
rect 25096 26404 25145 26432
rect 25096 26392 25102 26404
rect 25133 26401 25145 26404
rect 25179 26401 25191 26435
rect 25133 26395 25191 26401
rect 13446 26324 13452 26376
rect 13504 26364 13510 26376
rect 16224 26364 16252 26392
rect 13504 26336 16252 26364
rect 13504 26324 13510 26336
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 9398 26296 9404 26308
rect 8536 26268 9404 26296
rect 8536 26256 8542 26268
rect 9398 26256 9404 26268
rect 9456 26256 9462 26308
rect 11238 26296 11244 26308
rect 10626 26268 11244 26296
rect 11238 26256 11244 26268
rect 11296 26256 11302 26308
rect 14645 26299 14703 26305
rect 14645 26265 14657 26299
rect 14691 26296 14703 26299
rect 16025 26299 16083 26305
rect 14691 26268 15976 26296
rect 14691 26265 14703 26268
rect 14645 26259 14703 26265
rect 14737 26231 14795 26237
rect 14737 26197 14749 26231
rect 14783 26228 14795 26231
rect 14918 26228 14924 26240
rect 14783 26200 14924 26228
rect 14783 26197 14795 26200
rect 14737 26191 14795 26197
rect 14918 26188 14924 26200
rect 14976 26188 14982 26240
rect 15948 26228 15976 26268
rect 16025 26265 16037 26299
rect 16071 26296 16083 26299
rect 16390 26296 16396 26308
rect 16071 26268 16396 26296
rect 16071 26265 16083 26268
rect 16025 26259 16083 26265
rect 16390 26256 16396 26268
rect 16448 26256 16454 26308
rect 16960 26296 16988 26392
rect 18322 26324 18328 26376
rect 18380 26324 18386 26376
rect 19426 26324 19432 26376
rect 19484 26324 19490 26376
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 23290 26364 23296 26376
rect 23155 26336 23296 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 23290 26324 23296 26336
rect 23348 26324 23354 26376
rect 23842 26324 23848 26376
rect 23900 26324 23906 26376
rect 26050 26364 26056 26376
rect 23952 26336 26056 26364
rect 17310 26296 17316 26308
rect 16500 26268 17316 26296
rect 16500 26228 16528 26268
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 18340 26296 18368 26324
rect 20162 26296 20168 26308
rect 18340 26268 20168 26296
rect 20162 26256 20168 26268
rect 20220 26256 20226 26308
rect 22370 26256 22376 26308
rect 22428 26296 22434 26308
rect 23017 26299 23075 26305
rect 23017 26296 23029 26299
rect 22428 26268 23029 26296
rect 22428 26256 22434 26268
rect 23017 26265 23029 26268
rect 23063 26296 23075 26299
rect 23952 26296 23980 26336
rect 26050 26324 26056 26336
rect 26108 26324 26114 26376
rect 23063 26268 23980 26296
rect 25041 26299 25099 26305
rect 23063 26265 23075 26268
rect 23017 26259 23075 26265
rect 25041 26265 25053 26299
rect 25087 26296 25099 26299
rect 25130 26296 25136 26308
rect 25087 26268 25136 26296
rect 25087 26265 25099 26268
rect 25041 26259 25099 26265
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 15948 26200 16528 26228
rect 18233 26231 18291 26237
rect 18233 26197 18245 26231
rect 18279 26228 18291 26231
rect 18322 26228 18328 26240
rect 18279 26200 18328 26228
rect 18279 26197 18291 26200
rect 18233 26191 18291 26197
rect 18322 26188 18328 26200
rect 18380 26188 18386 26240
rect 24949 26231 25007 26237
rect 24949 26197 24961 26231
rect 24995 26228 25007 26231
rect 25866 26228 25872 26240
rect 24995 26200 25872 26228
rect 24995 26197 25007 26200
rect 24949 26191 25007 26197
rect 25866 26188 25872 26200
rect 25924 26188 25930 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 12437 26027 12495 26033
rect 12437 25993 12449 26027
rect 12483 26024 12495 26027
rect 12618 26024 12624 26036
rect 12483 25996 12624 26024
rect 12483 25993 12495 25996
rect 12437 25987 12495 25993
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 12897 26027 12955 26033
rect 12897 25993 12909 26027
rect 12943 26024 12955 26027
rect 16850 26024 16856 26036
rect 12943 25996 16856 26024
rect 12943 25993 12955 25996
rect 12897 25987 12955 25993
rect 16850 25984 16856 25996
rect 16908 25984 16914 26036
rect 18141 26027 18199 26033
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 18322 26024 18328 26036
rect 18187 25996 18328 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 19058 25984 19064 26036
rect 19116 26024 19122 26036
rect 22186 26024 22192 26036
rect 19116 25996 22192 26024
rect 19116 25984 19122 25996
rect 22186 25984 22192 25996
rect 22244 25984 22250 26036
rect 22462 25984 22468 26036
rect 22520 25984 22526 26036
rect 24762 26024 24768 26036
rect 23400 25996 24768 26024
rect 11422 25916 11428 25968
rect 11480 25956 11486 25968
rect 13909 25959 13967 25965
rect 13909 25956 13921 25959
rect 11480 25928 13921 25956
rect 11480 25916 11486 25928
rect 13909 25925 13921 25928
rect 13955 25925 13967 25959
rect 13909 25919 13967 25925
rect 15289 25959 15347 25965
rect 15289 25925 15301 25959
rect 15335 25956 15347 25959
rect 18233 25959 18291 25965
rect 15335 25928 16160 25956
rect 15335 25925 15347 25928
rect 15289 25919 15347 25925
rect 9950 25848 9956 25900
rect 10008 25888 10014 25900
rect 12529 25891 12587 25897
rect 12529 25888 12541 25891
rect 10008 25860 12541 25888
rect 10008 25848 10014 25860
rect 12529 25857 12541 25860
rect 12575 25857 12587 25891
rect 12529 25851 12587 25857
rect 13817 25891 13875 25897
rect 13817 25857 13829 25891
rect 13863 25888 13875 25891
rect 14642 25888 14648 25900
rect 13863 25860 14648 25888
rect 13863 25857 13875 25860
rect 13817 25851 13875 25857
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 15856 25888 15976 25892
rect 16025 25891 16083 25897
rect 16025 25888 16037 25891
rect 15243 25864 16037 25888
rect 15243 25860 15884 25864
rect 15948 25860 16037 25864
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 16025 25857 16037 25860
rect 16071 25857 16083 25891
rect 16132 25888 16160 25928
rect 18233 25925 18245 25959
rect 18279 25956 18291 25959
rect 18966 25956 18972 25968
rect 18279 25928 18972 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 18966 25916 18972 25928
rect 19024 25916 19030 25968
rect 22373 25959 22431 25965
rect 22373 25956 22385 25959
rect 22066 25928 22385 25956
rect 16132 25860 16712 25888
rect 16025 25851 16083 25857
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 12253 25823 12311 25829
rect 12253 25820 12265 25823
rect 11112 25792 12265 25820
rect 11112 25780 11118 25792
rect 12253 25789 12265 25792
rect 12299 25789 12311 25823
rect 12253 25783 12311 25789
rect 13354 25780 13360 25832
rect 13412 25820 13418 25832
rect 13633 25823 13691 25829
rect 13633 25820 13645 25823
rect 13412 25792 13645 25820
rect 13412 25780 13418 25792
rect 13633 25789 13645 25792
rect 13679 25789 13691 25823
rect 13633 25783 13691 25789
rect 15378 25780 15384 25832
rect 15436 25780 15442 25832
rect 16684 25820 16712 25860
rect 16850 25848 16856 25900
rect 16908 25848 16914 25900
rect 21450 25848 21456 25900
rect 21508 25888 21514 25900
rect 22066 25888 22094 25928
rect 22373 25925 22385 25928
rect 22419 25956 22431 25959
rect 23400 25956 23428 25996
rect 24762 25984 24768 25996
rect 24820 25984 24826 26036
rect 24854 25956 24860 25968
rect 22419 25928 23428 25956
rect 23492 25928 24860 25956
rect 22419 25925 22431 25928
rect 22373 25919 22431 25925
rect 23492 25897 23520 25928
rect 24854 25916 24860 25928
rect 24912 25916 24918 25968
rect 21508 25860 22094 25888
rect 23477 25891 23535 25897
rect 21508 25848 21514 25860
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23934 25848 23940 25900
rect 23992 25848 23998 25900
rect 17402 25820 17408 25832
rect 16684 25792 17408 25820
rect 17402 25780 17408 25792
rect 17460 25820 17466 25832
rect 17460 25792 17724 25820
rect 17460 25780 17466 25792
rect 14277 25755 14335 25761
rect 14277 25721 14289 25755
rect 14323 25752 14335 25755
rect 17586 25752 17592 25764
rect 14323 25724 15332 25752
rect 14323 25721 14335 25724
rect 14277 25715 14335 25721
rect 13814 25644 13820 25696
rect 13872 25684 13878 25696
rect 14829 25687 14887 25693
rect 14829 25684 14841 25687
rect 13872 25656 14841 25684
rect 13872 25644 13878 25656
rect 14829 25653 14841 25656
rect 14875 25653 14887 25687
rect 15304 25684 15332 25724
rect 16960 25724 17592 25752
rect 16960 25684 16988 25724
rect 17586 25712 17592 25724
rect 17644 25712 17650 25764
rect 17696 25752 17724 25792
rect 18414 25780 18420 25832
rect 18472 25780 18478 25832
rect 20898 25780 20904 25832
rect 20956 25820 20962 25832
rect 22557 25823 22615 25829
rect 20956 25792 22324 25820
rect 20956 25780 20962 25792
rect 22296 25752 22324 25792
rect 22557 25789 22569 25823
rect 22603 25789 22615 25823
rect 22557 25783 22615 25789
rect 22572 25752 22600 25783
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 25590 25752 25596 25764
rect 17696 25724 22232 25752
rect 22296 25724 22600 25752
rect 22664 25724 25596 25752
rect 15304 25656 16988 25684
rect 14829 25647 14887 25653
rect 17034 25644 17040 25696
rect 17092 25644 17098 25696
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 17773 25687 17831 25693
rect 17773 25684 17785 25687
rect 17460 25656 17785 25684
rect 17460 25644 17466 25656
rect 17773 25653 17785 25656
rect 17819 25653 17831 25687
rect 17773 25647 17831 25653
rect 18322 25644 18328 25696
rect 18380 25684 18386 25696
rect 19058 25684 19064 25696
rect 18380 25656 19064 25684
rect 18380 25644 18386 25656
rect 19058 25644 19064 25656
rect 19116 25644 19122 25696
rect 21450 25644 21456 25696
rect 21508 25684 21514 25696
rect 21545 25687 21603 25693
rect 21545 25684 21557 25687
rect 21508 25656 21557 25684
rect 21508 25644 21514 25656
rect 21545 25653 21557 25656
rect 21591 25653 21603 25687
rect 21545 25647 21603 25653
rect 22002 25644 22008 25696
rect 22060 25644 22066 25696
rect 22204 25684 22232 25724
rect 22664 25684 22692 25724
rect 25590 25712 25596 25724
rect 25648 25712 25654 25764
rect 22204 25656 22692 25684
rect 23293 25687 23351 25693
rect 23293 25653 23305 25687
rect 23339 25684 23351 25687
rect 23382 25684 23388 25696
rect 23339 25656 23388 25684
rect 23339 25653 23351 25656
rect 23293 25647 23351 25653
rect 23382 25644 23388 25656
rect 23440 25644 23446 25696
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 11698 25440 11704 25492
rect 11756 25480 11762 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 11756 25452 14289 25480
rect 11756 25440 11762 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 17129 25483 17187 25489
rect 17129 25449 17141 25483
rect 17175 25480 17187 25483
rect 21542 25480 21548 25492
rect 17175 25452 21548 25480
rect 17175 25449 17187 25452
rect 17129 25443 17187 25449
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 21729 25483 21787 25489
rect 21729 25449 21741 25483
rect 21775 25480 21787 25483
rect 23934 25480 23940 25492
rect 21775 25452 23940 25480
rect 21775 25449 21787 25452
rect 21729 25443 21787 25449
rect 23934 25440 23940 25452
rect 23992 25440 23998 25492
rect 24489 25483 24547 25489
rect 24489 25449 24501 25483
rect 24535 25480 24547 25483
rect 24854 25480 24860 25492
rect 24535 25452 24860 25480
rect 24535 25449 24547 25452
rect 24489 25443 24547 25449
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 25774 25480 25780 25492
rect 25648 25452 25780 25480
rect 25648 25440 25654 25452
rect 25774 25440 25780 25452
rect 25832 25440 25838 25492
rect 14642 25372 14648 25424
rect 14700 25412 14706 25424
rect 15194 25412 15200 25424
rect 14700 25384 15200 25412
rect 14700 25372 14706 25384
rect 15194 25372 15200 25384
rect 15252 25372 15258 25424
rect 18141 25415 18199 25421
rect 18141 25412 18153 25415
rect 16868 25384 18153 25412
rect 14734 25304 14740 25356
rect 14792 25344 14798 25356
rect 14829 25347 14887 25353
rect 14829 25344 14841 25347
rect 14792 25316 14841 25344
rect 14792 25304 14798 25316
rect 14829 25313 14841 25316
rect 14875 25313 14887 25347
rect 14829 25307 14887 25313
rect 16301 25347 16359 25353
rect 16301 25313 16313 25347
rect 16347 25313 16359 25347
rect 16301 25307 16359 25313
rect 11238 25236 11244 25288
rect 11296 25236 11302 25288
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25245 12679 25279
rect 12621 25239 12679 25245
rect 12345 25211 12403 25217
rect 12345 25177 12357 25211
rect 12391 25177 12403 25211
rect 12636 25208 12664 25239
rect 12802 25236 12808 25288
rect 12860 25276 12866 25288
rect 16316 25276 16344 25307
rect 12860 25248 16344 25276
rect 12860 25236 12866 25248
rect 14826 25208 14832 25220
rect 12636 25180 14832 25208
rect 12345 25171 12403 25177
rect 9674 25100 9680 25152
rect 9732 25140 9738 25152
rect 10778 25140 10784 25152
rect 9732 25112 10784 25140
rect 9732 25100 9738 25112
rect 10778 25100 10784 25112
rect 10836 25140 10842 25152
rect 10873 25143 10931 25149
rect 10873 25140 10885 25143
rect 10836 25112 10885 25140
rect 10836 25100 10842 25112
rect 10873 25109 10885 25112
rect 10919 25109 10931 25143
rect 12360 25140 12388 25171
rect 14826 25168 14832 25180
rect 14884 25168 14890 25220
rect 15838 25208 15844 25220
rect 15212 25180 15844 25208
rect 12894 25140 12900 25152
rect 12360 25112 12900 25140
rect 10873 25103 10931 25109
rect 12894 25100 12900 25112
rect 12952 25100 12958 25152
rect 12986 25100 12992 25152
rect 13044 25100 13050 25152
rect 14642 25100 14648 25152
rect 14700 25100 14706 25152
rect 14737 25143 14795 25149
rect 14737 25109 14749 25143
rect 14783 25140 14795 25143
rect 15212 25140 15240 25180
rect 15838 25168 15844 25180
rect 15896 25168 15902 25220
rect 16117 25211 16175 25217
rect 16117 25177 16129 25211
rect 16163 25208 16175 25211
rect 16868 25208 16896 25384
rect 18141 25381 18153 25384
rect 18187 25412 18199 25415
rect 18598 25412 18604 25424
rect 18187 25384 18604 25412
rect 18187 25381 18199 25384
rect 18141 25375 18199 25381
rect 18598 25372 18604 25384
rect 18656 25412 18662 25424
rect 19337 25415 19395 25421
rect 19337 25412 19349 25415
rect 18656 25384 19349 25412
rect 18656 25372 18662 25384
rect 19337 25381 19349 25384
rect 19383 25412 19395 25415
rect 19886 25412 19892 25424
rect 19383 25384 19892 25412
rect 19383 25381 19395 25384
rect 19337 25375 19395 25381
rect 19886 25372 19892 25384
rect 19944 25372 19950 25424
rect 20346 25372 20352 25424
rect 20404 25372 20410 25424
rect 20993 25415 21051 25421
rect 20993 25412 21005 25415
rect 20916 25384 21005 25412
rect 17034 25304 17040 25356
rect 17092 25344 17098 25356
rect 17092 25316 20852 25344
rect 17092 25304 17098 25316
rect 16942 25236 16948 25288
rect 17000 25236 17006 25288
rect 17586 25236 17592 25288
rect 17644 25236 17650 25288
rect 18322 25276 18328 25288
rect 17696 25248 18328 25276
rect 16163 25180 16896 25208
rect 16163 25177 16175 25180
rect 16117 25171 16175 25177
rect 14783 25112 15240 25140
rect 14783 25109 14795 25112
rect 14737 25103 14795 25109
rect 15286 25100 15292 25152
rect 15344 25100 15350 25152
rect 15746 25100 15752 25152
rect 15804 25100 15810 25152
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16298 25140 16304 25152
rect 16255 25112 16304 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 16298 25100 16304 25112
rect 16356 25140 16362 25152
rect 17696 25140 17724 25248
rect 18322 25236 18328 25248
rect 18380 25236 18386 25288
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20346 25276 20352 25288
rect 19935 25248 20352 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20346 25236 20352 25248
rect 20404 25236 20410 25288
rect 20824 25285 20852 25316
rect 20809 25279 20867 25285
rect 20809 25245 20821 25279
rect 20855 25245 20867 25279
rect 20809 25239 20867 25245
rect 17788 25180 19334 25208
rect 17788 25149 17816 25180
rect 16356 25112 17724 25140
rect 17773 25143 17831 25149
rect 16356 25100 16362 25112
rect 17773 25109 17785 25143
rect 17819 25109 17831 25143
rect 17773 25103 17831 25109
rect 18322 25100 18328 25152
rect 18380 25100 18386 25152
rect 18506 25100 18512 25152
rect 18564 25140 18570 25152
rect 18693 25143 18751 25149
rect 18693 25140 18705 25143
rect 18564 25112 18705 25140
rect 18564 25100 18570 25112
rect 18693 25109 18705 25112
rect 18739 25109 18751 25143
rect 19306 25140 19334 25180
rect 19702 25168 19708 25220
rect 19760 25168 19766 25220
rect 20916 25208 20944 25384
rect 20993 25381 21005 25384
rect 21039 25381 21051 25415
rect 20993 25375 21051 25381
rect 23842 25372 23848 25424
rect 23900 25412 23906 25424
rect 24581 25415 24639 25421
rect 24581 25412 24593 25415
rect 23900 25384 24593 25412
rect 23900 25372 23906 25384
rect 24581 25381 24593 25384
rect 24627 25381 24639 25415
rect 24581 25375 24639 25381
rect 24670 25372 24676 25424
rect 24728 25412 24734 25424
rect 25133 25415 25191 25421
rect 25133 25412 25145 25415
rect 24728 25384 25145 25412
rect 24728 25372 24734 25384
rect 25133 25381 25145 25384
rect 25179 25381 25191 25415
rect 25133 25375 25191 25381
rect 21542 25236 21548 25288
rect 21600 25236 21606 25288
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22664 25208 22692 25239
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 20916 25180 22692 25208
rect 23842 25168 23848 25220
rect 23900 25168 23906 25220
rect 22186 25140 22192 25152
rect 19306 25112 22192 25140
rect 18693 25103 18751 25109
rect 22186 25100 22192 25112
rect 22244 25100 22250 25152
rect 24857 25143 24915 25149
rect 24857 25109 24869 25143
rect 24903 25140 24915 25143
rect 25498 25140 25504 25152
rect 24903 25112 25504 25140
rect 24903 25109 24915 25112
rect 24857 25103 24915 25109
rect 25498 25100 25504 25112
rect 25556 25140 25562 25152
rect 25866 25140 25872 25152
rect 25556 25112 25872 25140
rect 25556 25100 25562 25112
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 10502 24896 10508 24948
rect 10560 24936 10566 24948
rect 15286 24936 15292 24948
rect 10560 24908 15292 24936
rect 10560 24896 10566 24908
rect 15286 24896 15292 24908
rect 15344 24896 15350 24948
rect 17218 24896 17224 24948
rect 17276 24896 17282 24948
rect 18417 24939 18475 24945
rect 18417 24905 18429 24939
rect 18463 24936 18475 24939
rect 19886 24936 19892 24948
rect 18463 24908 19892 24936
rect 18463 24905 18475 24908
rect 18417 24899 18475 24905
rect 19886 24896 19892 24908
rect 19944 24896 19950 24948
rect 11790 24828 11796 24880
rect 11848 24868 11854 24880
rect 12069 24871 12127 24877
rect 12069 24868 12081 24871
rect 11848 24840 12081 24868
rect 11848 24828 11854 24840
rect 12069 24837 12081 24840
rect 12115 24837 12127 24871
rect 12069 24831 12127 24837
rect 12710 24828 12716 24880
rect 12768 24868 12774 24880
rect 12986 24868 12992 24880
rect 12768 24840 12992 24868
rect 12768 24828 12774 24840
rect 12986 24828 12992 24840
rect 13044 24868 13050 24880
rect 17236 24868 17264 24896
rect 18598 24868 18604 24880
rect 13044 24840 13294 24868
rect 17236 24840 18604 24868
rect 13044 24828 13050 24840
rect 18598 24828 18604 24840
rect 18656 24868 18662 24880
rect 18656 24840 19104 24868
rect 18656 24828 18662 24840
rect 9122 24760 9128 24812
rect 9180 24800 9186 24812
rect 9180 24772 9798 24800
rect 9180 24760 9186 24772
rect 11974 24760 11980 24812
rect 12032 24760 12038 24812
rect 14737 24803 14795 24809
rect 14737 24769 14749 24803
rect 14783 24800 14795 24803
rect 14826 24800 14832 24812
rect 14783 24772 14832 24800
rect 14783 24769 14795 24772
rect 14737 24763 14795 24769
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 15194 24760 15200 24812
rect 15252 24760 15258 24812
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24800 15439 24803
rect 15838 24800 15844 24812
rect 15427 24772 15844 24800
rect 15427 24769 15439 24772
rect 15381 24763 15439 24769
rect 15838 24760 15844 24772
rect 15896 24800 15902 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 15896 24772 17325 24800
rect 15896 24760 15902 24772
rect 17313 24769 17325 24772
rect 17359 24800 17371 24803
rect 17359 24772 17908 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 10873 24735 10931 24741
rect 10873 24701 10885 24735
rect 10919 24732 10931 24735
rect 10919 24704 11100 24732
rect 10919 24701 10931 24704
rect 10873 24695 10931 24701
rect 11072 24608 11100 24704
rect 11146 24692 11152 24744
rect 11204 24692 11210 24744
rect 11885 24735 11943 24741
rect 11885 24701 11897 24735
rect 11931 24732 11943 24735
rect 12066 24732 12072 24744
rect 11931 24704 12072 24732
rect 11931 24701 11943 24704
rect 11885 24695 11943 24701
rect 12066 24692 12072 24704
rect 12124 24692 12130 24744
rect 12894 24692 12900 24744
rect 12952 24732 12958 24744
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12952 24704 13001 24732
rect 12952 24692 12958 24704
rect 12989 24701 13001 24704
rect 13035 24732 13047 24735
rect 13446 24732 13452 24744
rect 13035 24704 13452 24732
rect 13035 24701 13047 24704
rect 12989 24695 13047 24701
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 13722 24692 13728 24744
rect 13780 24732 13786 24744
rect 14461 24735 14519 24741
rect 14461 24732 14473 24735
rect 13780 24704 14473 24732
rect 13780 24692 13786 24704
rect 14461 24701 14473 24704
rect 14507 24701 14519 24735
rect 16942 24732 16948 24744
rect 14461 24695 14519 24701
rect 14660 24704 16948 24732
rect 12437 24667 12495 24673
rect 12437 24633 12449 24667
rect 12483 24664 12495 24667
rect 12483 24636 13492 24664
rect 12483 24633 12495 24636
rect 12437 24627 12495 24633
rect 9398 24556 9404 24608
rect 9456 24556 9462 24608
rect 11054 24556 11060 24608
rect 11112 24556 11118 24608
rect 13464 24596 13492 24636
rect 14660 24596 14688 24704
rect 16942 24692 16948 24704
rect 17000 24692 17006 24744
rect 17034 24692 17040 24744
rect 17092 24732 17098 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 17092 24704 17417 24732
rect 17092 24692 17098 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17880 24732 17908 24772
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 19076 24809 19104 24840
rect 20254 24828 20260 24880
rect 20312 24868 20318 24880
rect 22465 24871 22523 24877
rect 20312 24840 20470 24868
rect 20312 24828 20318 24840
rect 22465 24837 22477 24871
rect 22511 24868 22523 24871
rect 24118 24868 24124 24880
rect 22511 24840 24124 24868
rect 22511 24837 22523 24840
rect 22465 24831 22523 24837
rect 24118 24828 24124 24840
rect 24176 24828 24182 24880
rect 18509 24803 18567 24809
rect 18509 24800 18521 24803
rect 18380 24772 18521 24800
rect 18380 24760 18386 24772
rect 18509 24769 18521 24772
rect 18555 24800 18567 24803
rect 19061 24803 19119 24809
rect 18555 24772 18736 24800
rect 18555 24769 18567 24772
rect 18509 24763 18567 24769
rect 18414 24732 18420 24744
rect 17880 24704 18420 24732
rect 17405 24695 17463 24701
rect 18414 24692 18420 24704
rect 18472 24692 18478 24744
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24701 18659 24735
rect 18601 24695 18659 24701
rect 15378 24624 15384 24676
rect 15436 24664 15442 24676
rect 16853 24667 16911 24673
rect 16853 24664 16865 24667
rect 15436 24636 16865 24664
rect 15436 24624 15442 24636
rect 16853 24633 16865 24636
rect 16899 24633 16911 24667
rect 18616 24664 18644 24695
rect 16853 24627 16911 24633
rect 16960 24636 18644 24664
rect 18708 24664 18736 24772
rect 19061 24769 19073 24803
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 22646 24800 22652 24812
rect 22603 24772 22652 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 22646 24760 22652 24772
rect 22704 24760 22710 24812
rect 24946 24760 24952 24812
rect 25004 24760 25010 24812
rect 19150 24692 19156 24744
rect 19208 24732 19214 24744
rect 19426 24732 19432 24744
rect 19208 24704 19432 24732
rect 19208 24692 19214 24704
rect 19426 24692 19432 24704
rect 19484 24732 19490 24744
rect 19705 24735 19763 24741
rect 19705 24732 19717 24735
rect 19484 24704 19717 24732
rect 19484 24692 19490 24704
rect 19705 24701 19717 24704
rect 19751 24701 19763 24735
rect 19705 24695 19763 24701
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20070 24732 20076 24744
rect 20027 24704 20076 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 22278 24732 22284 24744
rect 21499 24704 22284 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 22278 24692 22284 24704
rect 22336 24692 22342 24744
rect 22738 24692 22744 24744
rect 22796 24692 22802 24744
rect 23290 24692 23296 24744
rect 23348 24732 23354 24744
rect 23566 24732 23572 24744
rect 23348 24704 23572 24732
rect 23348 24692 23354 24704
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 25038 24732 25044 24744
rect 23891 24704 25044 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 25317 24735 25375 24741
rect 25317 24701 25329 24735
rect 25363 24732 25375 24735
rect 25406 24732 25412 24744
rect 25363 24704 25412 24732
rect 25363 24701 25375 24704
rect 25317 24695 25375 24701
rect 25406 24692 25412 24704
rect 25464 24692 25470 24744
rect 18708 24636 19748 24664
rect 13464 24568 14688 24596
rect 15470 24556 15476 24608
rect 15528 24556 15534 24608
rect 16482 24556 16488 24608
rect 16540 24596 16546 24608
rect 16960 24596 16988 24636
rect 19720 24608 19748 24636
rect 21542 24624 21548 24676
rect 21600 24664 21606 24676
rect 23201 24667 23259 24673
rect 23201 24664 23213 24667
rect 21600 24636 23213 24664
rect 21600 24624 21606 24636
rect 23201 24633 23213 24636
rect 23247 24633 23259 24667
rect 23201 24627 23259 24633
rect 16540 24568 16988 24596
rect 18049 24599 18107 24605
rect 16540 24556 16546 24568
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18322 24596 18328 24608
rect 18095 24568 18328 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 18414 24556 18420 24608
rect 18472 24596 18478 24608
rect 19337 24599 19395 24605
rect 19337 24596 19349 24599
rect 18472 24568 19349 24596
rect 18472 24556 18478 24568
rect 19337 24565 19349 24568
rect 19383 24565 19395 24599
rect 19337 24559 19395 24565
rect 19702 24556 19708 24608
rect 19760 24556 19766 24608
rect 21358 24556 21364 24608
rect 21416 24596 21422 24608
rect 22097 24599 22155 24605
rect 22097 24596 22109 24599
rect 21416 24568 22109 24596
rect 21416 24556 21422 24568
rect 22097 24565 22109 24568
rect 22143 24565 22155 24599
rect 22097 24559 22155 24565
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 9398 24352 9404 24404
rect 9456 24392 9462 24404
rect 9582 24392 9588 24404
rect 9456 24364 9588 24392
rect 9456 24352 9462 24364
rect 9582 24352 9588 24364
rect 9640 24392 9646 24404
rect 9640 24364 13676 24392
rect 9640 24352 9646 24364
rect 13648 24324 13676 24364
rect 13722 24352 13728 24404
rect 13780 24352 13786 24404
rect 21634 24392 21640 24404
rect 19076 24364 21640 24392
rect 14734 24324 14740 24336
rect 13648 24296 14740 24324
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 18141 24327 18199 24333
rect 18141 24293 18153 24327
rect 18187 24324 18199 24327
rect 18874 24324 18880 24336
rect 18187 24296 18880 24324
rect 18187 24293 18199 24296
rect 18141 24287 18199 24293
rect 18874 24284 18880 24296
rect 18932 24284 18938 24336
rect 11146 24216 11152 24268
rect 11204 24256 11210 24268
rect 11977 24259 12035 24265
rect 11977 24256 11989 24259
rect 11204 24228 11989 24256
rect 11204 24216 11210 24228
rect 11977 24225 11989 24228
rect 12023 24256 12035 24259
rect 12342 24256 12348 24268
rect 12023 24228 12348 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 12710 24216 12716 24268
rect 12768 24256 12774 24268
rect 14093 24259 14151 24265
rect 14093 24256 14105 24259
rect 12768 24228 14105 24256
rect 12768 24216 12774 24228
rect 14093 24225 14105 24228
rect 14139 24256 14151 24259
rect 15470 24256 15476 24268
rect 14139 24228 15476 24256
rect 14139 24225 14151 24228
rect 14093 24219 14151 24225
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 18690 24216 18696 24268
rect 18748 24216 18754 24268
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 7892 24160 9137 24188
rect 7892 24148 7898 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 19076 24188 19104 24364
rect 21634 24352 21640 24364
rect 21692 24352 21698 24404
rect 24029 24395 24087 24401
rect 24029 24361 24041 24395
rect 24075 24392 24087 24395
rect 24946 24392 24952 24404
rect 24075 24364 24952 24392
rect 24075 24361 24087 24364
rect 24029 24355 24087 24361
rect 24946 24352 24952 24364
rect 25004 24392 25010 24404
rect 25130 24392 25136 24404
rect 25004 24364 25136 24392
rect 25004 24352 25010 24364
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 25314 24352 25320 24404
rect 25372 24392 25378 24404
rect 25409 24395 25467 24401
rect 25409 24392 25421 24395
rect 25372 24364 25421 24392
rect 25372 24352 25378 24364
rect 25409 24361 25421 24364
rect 25455 24361 25467 24395
rect 25409 24355 25467 24361
rect 23290 24284 23296 24336
rect 23348 24284 23354 24336
rect 19150 24216 19156 24268
rect 19208 24256 19214 24268
rect 21177 24259 21235 24265
rect 21177 24256 21189 24259
rect 19208 24228 21189 24256
rect 19208 24216 19214 24228
rect 21177 24225 21189 24228
rect 21223 24225 21235 24259
rect 21177 24219 21235 24225
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 23308 24256 23336 24284
rect 21959 24228 23336 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24176 24228 24593 24256
rect 24176 24216 24182 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 18647 24160 19104 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 9401 24123 9459 24129
rect 9401 24089 9413 24123
rect 9447 24120 9459 24123
rect 9490 24120 9496 24132
rect 9447 24092 9496 24120
rect 9447 24089 9459 24092
rect 9401 24083 9459 24089
rect 9490 24080 9496 24092
rect 9548 24080 9554 24132
rect 11238 24120 11244 24132
rect 9784 24092 9890 24120
rect 10704 24092 11244 24120
rect 8386 24012 8392 24064
rect 8444 24052 8450 24064
rect 9122 24052 9128 24064
rect 8444 24024 9128 24052
rect 8444 24012 8450 24024
rect 9122 24012 9128 24024
rect 9180 24052 9186 24064
rect 9784 24052 9812 24092
rect 10704 24052 10732 24092
rect 11238 24080 11244 24092
rect 11296 24120 11302 24132
rect 11425 24123 11483 24129
rect 11425 24120 11437 24123
rect 11296 24092 11437 24120
rect 11296 24080 11302 24092
rect 11425 24089 11437 24092
rect 11471 24089 11483 24123
rect 11425 24083 11483 24089
rect 11514 24080 11520 24132
rect 11572 24120 11578 24132
rect 12253 24123 12311 24129
rect 12253 24120 12265 24123
rect 11572 24092 12265 24120
rect 11572 24080 11578 24092
rect 12253 24089 12265 24092
rect 12299 24120 12311 24123
rect 12526 24120 12532 24132
rect 12299 24092 12532 24120
rect 12299 24089 12311 24092
rect 12253 24083 12311 24089
rect 12526 24080 12532 24092
rect 12584 24080 12590 24132
rect 12710 24080 12716 24132
rect 12768 24080 12774 24132
rect 17681 24123 17739 24129
rect 17681 24089 17693 24123
rect 17727 24120 17739 24123
rect 18966 24120 18972 24132
rect 17727 24092 18972 24120
rect 17727 24089 17739 24092
rect 17681 24083 17739 24089
rect 18966 24080 18972 24092
rect 19024 24080 19030 24132
rect 20346 24080 20352 24132
rect 20404 24080 20410 24132
rect 20438 24080 20444 24132
rect 20496 24120 20502 24132
rect 20496 24092 20852 24120
rect 20496 24080 20502 24092
rect 9180 24024 10732 24052
rect 10873 24055 10931 24061
rect 9180 24012 9186 24024
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11146 24052 11152 24064
rect 10919 24024 11152 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 16393 24055 16451 24061
rect 16393 24021 16405 24055
rect 16439 24052 16451 24055
rect 16666 24052 16672 24064
rect 16439 24024 16672 24052
rect 16439 24021 16451 24024
rect 16393 24015 16451 24021
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 16758 24012 16764 24064
rect 16816 24052 16822 24064
rect 18506 24052 18512 24064
rect 16816 24024 18512 24052
rect 16816 24012 16822 24024
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 20070 24052 20076 24064
rect 19475 24024 20076 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 20070 24012 20076 24024
rect 20128 24012 20134 24064
rect 20824 24052 20852 24092
rect 20898 24080 20904 24132
rect 20956 24080 20962 24132
rect 22189 24123 22247 24129
rect 22189 24089 22201 24123
rect 22235 24120 22247 24123
rect 22278 24120 22284 24132
rect 22235 24092 22284 24120
rect 22235 24089 22247 24092
rect 22189 24083 22247 24089
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 22388 24092 22678 24120
rect 21542 24052 21548 24064
rect 20824 24024 21548 24052
rect 21542 24012 21548 24024
rect 21600 24052 21606 24064
rect 22388 24052 22416 24092
rect 21600 24024 22416 24052
rect 21600 24012 21606 24024
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23532 24024 23673 24052
rect 23532 24012 23538 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 10045 23851 10103 23857
rect 10045 23848 10057 23851
rect 8680 23820 10057 23848
rect 8386 23740 8392 23792
rect 8444 23780 8450 23792
rect 8680 23780 8708 23820
rect 10045 23817 10057 23820
rect 10091 23817 10103 23851
rect 10045 23811 10103 23817
rect 10410 23808 10416 23860
rect 10468 23808 10474 23860
rect 13354 23808 13360 23860
rect 13412 23848 13418 23860
rect 14737 23851 14795 23857
rect 13412 23820 13860 23848
rect 13412 23808 13418 23820
rect 8444 23752 8786 23780
rect 8444 23740 8450 23752
rect 13630 23740 13636 23792
rect 13688 23740 13694 23792
rect 13722 23740 13728 23792
rect 13780 23740 13786 23792
rect 13832 23780 13860 23820
rect 14737 23817 14749 23851
rect 14783 23848 14795 23851
rect 15010 23848 15016 23860
rect 14783 23820 15016 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 15010 23808 15016 23820
rect 15068 23808 15074 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 16816 23820 17233 23848
rect 16816 23808 16822 23820
rect 17221 23817 17233 23820
rect 17267 23817 17279 23851
rect 17221 23811 17279 23817
rect 17313 23851 17371 23857
rect 17313 23817 17325 23851
rect 17359 23848 17371 23851
rect 17494 23848 17500 23860
rect 17359 23820 17500 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 17494 23808 17500 23820
rect 17552 23848 17558 23860
rect 17862 23848 17868 23860
rect 17552 23820 17868 23848
rect 17552 23808 17558 23820
rect 17862 23808 17868 23820
rect 17920 23848 17926 23860
rect 18693 23851 18751 23857
rect 18693 23848 18705 23851
rect 17920 23820 18705 23848
rect 17920 23808 17926 23820
rect 18693 23817 18705 23820
rect 18739 23817 18751 23851
rect 18693 23811 18751 23817
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23817 20039 23851
rect 19981 23811 20039 23817
rect 20901 23851 20959 23857
rect 20901 23817 20913 23851
rect 20947 23848 20959 23851
rect 21910 23848 21916 23860
rect 20947 23820 21916 23848
rect 20947 23817 20959 23820
rect 20901 23811 20959 23817
rect 14829 23783 14887 23789
rect 14829 23780 14841 23783
rect 13832 23752 14841 23780
rect 14829 23749 14841 23752
rect 14875 23749 14887 23783
rect 14829 23743 14887 23749
rect 14918 23740 14924 23792
rect 14976 23780 14982 23792
rect 14976 23752 17448 23780
rect 14976 23740 14982 23752
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23712 10839 23715
rect 13538 23712 13544 23724
rect 10827 23684 13544 23712
rect 10827 23681 10839 23684
rect 10781 23675 10839 23681
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13740 23712 13768 23740
rect 17034 23712 17040 23724
rect 13740 23684 14596 23712
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 8021 23647 8079 23653
rect 8021 23644 8033 23647
rect 7892 23616 8033 23644
rect 7892 23604 7898 23616
rect 8021 23613 8033 23616
rect 8067 23613 8079 23647
rect 8021 23607 8079 23613
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23644 8355 23647
rect 10502 23644 10508 23656
rect 8343 23616 10508 23644
rect 8343 23613 8355 23616
rect 8297 23607 8355 23613
rect 10502 23604 10508 23616
rect 10560 23604 10566 23656
rect 10870 23604 10876 23656
rect 10928 23604 10934 23656
rect 10962 23604 10968 23656
rect 11020 23604 11026 23656
rect 13446 23604 13452 23656
rect 13504 23644 13510 23656
rect 14568 23653 14596 23684
rect 14660 23684 17040 23712
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 13504 23616 13737 23644
rect 13504 23604 13510 23616
rect 13725 23613 13737 23616
rect 13771 23613 13783 23647
rect 13725 23607 13783 23613
rect 13817 23647 13875 23653
rect 13817 23613 13829 23647
rect 13863 23613 13875 23647
rect 13817 23607 13875 23613
rect 14553 23647 14611 23653
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 9769 23579 9827 23585
rect 9769 23545 9781 23579
rect 9815 23576 9827 23579
rect 10980 23576 11008 23604
rect 13832 23576 13860 23607
rect 9815 23548 11008 23576
rect 12406 23548 13860 23576
rect 9815 23545 9827 23548
rect 9769 23539 9827 23545
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 12406 23508 12434 23548
rect 10836 23480 12434 23508
rect 10836 23468 10842 23480
rect 12526 23468 12532 23520
rect 12584 23508 12590 23520
rect 13265 23511 13323 23517
rect 13265 23508 13277 23511
rect 12584 23480 13277 23508
rect 12584 23468 12590 23480
rect 13265 23477 13277 23480
rect 13311 23477 13323 23511
rect 13265 23471 13323 23477
rect 13538 23468 13544 23520
rect 13596 23508 13602 23520
rect 14660 23508 14688 23684
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 15654 23604 15660 23656
rect 15712 23604 15718 23656
rect 17420 23653 17448 23752
rect 18506 23740 18512 23792
rect 18564 23780 18570 23792
rect 19242 23780 19248 23792
rect 18564 23752 19248 23780
rect 18564 23740 18570 23752
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 19996 23780 20024 23811
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 22925 23851 22983 23857
rect 22925 23817 22937 23851
rect 22971 23848 22983 23851
rect 24949 23851 25007 23857
rect 22971 23820 24808 23848
rect 22971 23817 22983 23820
rect 22925 23811 22983 23817
rect 20254 23780 20260 23792
rect 19444 23752 19748 23780
rect 19996 23752 20260 23780
rect 18049 23715 18107 23721
rect 18049 23681 18061 23715
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 15197 23579 15255 23585
rect 15197 23545 15209 23579
rect 15243 23576 15255 23579
rect 18064 23576 18092 23675
rect 19444 23653 19472 23752
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19720 23712 19748 23752
rect 20254 23740 20260 23752
rect 20312 23740 20318 23792
rect 20714 23740 20720 23792
rect 20772 23780 20778 23792
rect 20772 23752 21036 23780
rect 20772 23740 20778 23752
rect 19720 23684 20116 23712
rect 19429 23647 19487 23653
rect 19429 23613 19441 23647
rect 19475 23613 19487 23647
rect 19429 23607 19487 23613
rect 19521 23647 19579 23653
rect 19521 23613 19533 23647
rect 19567 23644 19579 23647
rect 19978 23644 19984 23656
rect 19567 23616 19984 23644
rect 19567 23613 19579 23616
rect 19521 23607 19579 23613
rect 19978 23604 19984 23616
rect 20036 23604 20042 23656
rect 20088 23644 20116 23684
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 20898 23644 20904 23656
rect 20088 23616 20904 23644
rect 20898 23604 20904 23616
rect 20956 23604 20962 23656
rect 21008 23653 21036 23752
rect 21542 23740 21548 23792
rect 21600 23780 21606 23792
rect 22940 23780 22968 23811
rect 24780 23780 24808 23820
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25038 23848 25044 23860
rect 24995 23820 25044 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25038 23808 25044 23820
rect 25096 23808 25102 23860
rect 25130 23780 25136 23792
rect 21600 23752 22968 23780
rect 24702 23752 25136 23780
rect 21600 23740 21606 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 22186 23672 22192 23724
rect 22244 23672 22250 23724
rect 20993 23647 21051 23653
rect 20993 23613 21005 23647
rect 21039 23613 21051 23647
rect 20993 23607 21051 23613
rect 23198 23604 23204 23656
rect 23256 23604 23262 23656
rect 23474 23604 23480 23656
rect 23532 23604 23538 23656
rect 15243 23548 18092 23576
rect 18233 23579 18291 23585
rect 15243 23545 15255 23548
rect 15197 23539 15255 23545
rect 18233 23545 18245 23579
rect 18279 23576 18291 23579
rect 18279 23548 19472 23576
rect 18279 23545 18291 23548
rect 18233 23539 18291 23545
rect 13596 23480 14688 23508
rect 16853 23511 16911 23517
rect 13596 23468 13602 23480
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 17126 23508 17132 23520
rect 16899 23480 17132 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 17126 23468 17132 23480
rect 17184 23468 17190 23520
rect 17310 23468 17316 23520
rect 17368 23508 17374 23520
rect 17494 23508 17500 23520
rect 17368 23480 17500 23508
rect 17368 23468 17374 23480
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 18138 23468 18144 23520
rect 18196 23508 18202 23520
rect 18414 23508 18420 23520
rect 18196 23480 18420 23508
rect 18196 23468 18202 23480
rect 18414 23468 18420 23480
rect 18472 23468 18478 23520
rect 18966 23468 18972 23520
rect 19024 23468 19030 23520
rect 19444 23508 19472 23548
rect 19794 23536 19800 23588
rect 19852 23576 19858 23588
rect 20441 23579 20499 23585
rect 20441 23576 20453 23579
rect 19852 23548 20453 23576
rect 19852 23536 19858 23548
rect 20441 23545 20453 23548
rect 20487 23545 20499 23579
rect 20441 23539 20499 23545
rect 22373 23579 22431 23585
rect 22373 23545 22385 23579
rect 22419 23576 22431 23579
rect 22419 23548 23152 23576
rect 22419 23545 22431 23548
rect 22373 23539 22431 23545
rect 21910 23508 21916 23520
rect 19444 23480 21916 23508
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 23124 23508 23152 23548
rect 23934 23508 23940 23520
rect 23124 23480 23940 23508
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 25130 23468 25136 23520
rect 25188 23508 25194 23520
rect 25225 23511 25283 23517
rect 25225 23508 25237 23511
rect 25188 23480 25237 23508
rect 25188 23468 25194 23480
rect 25225 23477 25237 23480
rect 25271 23508 25283 23511
rect 25498 23508 25504 23520
rect 25271 23480 25504 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 25498 23468 25504 23480
rect 25556 23468 25562 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9214 23304 9220 23316
rect 9171 23276 9220 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 10229 23307 10287 23313
rect 10229 23273 10241 23307
rect 10275 23304 10287 23307
rect 10502 23304 10508 23316
rect 10275 23276 10508 23304
rect 10275 23273 10287 23276
rect 10229 23267 10287 23273
rect 10502 23264 10508 23276
rect 10560 23264 10566 23316
rect 11054 23264 11060 23316
rect 11112 23304 11118 23316
rect 11330 23304 11336 23316
rect 11112 23276 11336 23304
rect 11112 23264 11118 23276
rect 11330 23264 11336 23276
rect 11388 23264 11394 23316
rect 11882 23264 11888 23316
rect 11940 23304 11946 23316
rect 14369 23307 14427 23313
rect 14369 23304 14381 23307
rect 11940 23276 14381 23304
rect 11940 23264 11946 23276
rect 14369 23273 14381 23276
rect 14415 23273 14427 23307
rect 14369 23267 14427 23273
rect 15841 23307 15899 23313
rect 15841 23273 15853 23307
rect 15887 23304 15899 23307
rect 17310 23304 17316 23316
rect 15887 23276 17316 23304
rect 15887 23273 15899 23276
rect 15841 23267 15899 23273
rect 8202 23196 8208 23248
rect 8260 23236 8266 23248
rect 8260 23208 11836 23236
rect 8260 23196 8266 23208
rect 8662 23128 8668 23180
rect 8720 23168 8726 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 8720 23140 9689 23168
rect 8720 23128 8726 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 11698 23128 11704 23180
rect 11756 23128 11762 23180
rect 11808 23177 11836 23208
rect 11793 23171 11851 23177
rect 11793 23137 11805 23171
rect 11839 23137 11851 23171
rect 11793 23131 11851 23137
rect 12986 23128 12992 23180
rect 13044 23168 13050 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13044 23140 13553 23168
rect 13044 23128 13050 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 14384 23168 14412 23267
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 14384 23140 15301 23168
rect 13541 23131 13599 23137
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 11606 23060 11612 23112
rect 11664 23060 11670 23112
rect 13449 23103 13507 23109
rect 13449 23069 13461 23103
rect 13495 23100 13507 23103
rect 14185 23103 14243 23109
rect 14185 23100 14197 23103
rect 13495 23072 14197 23100
rect 13495 23069 13507 23072
rect 13449 23063 13507 23069
rect 14185 23069 14197 23072
rect 14231 23100 14243 23103
rect 15105 23103 15163 23109
rect 14231 23072 15056 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 9493 23035 9551 23041
rect 9493 23001 9505 23035
rect 9539 23032 9551 23035
rect 10410 23032 10416 23044
rect 9539 23004 10416 23032
rect 9539 23001 9551 23004
rect 9493 22995 9551 23001
rect 10410 22992 10416 23004
rect 10468 22992 10474 23044
rect 11330 22992 11336 23044
rect 11388 23032 11394 23044
rect 15028 23032 15056 23072
rect 15105 23069 15117 23103
rect 15151 23100 15163 23103
rect 15654 23100 15660 23112
rect 15151 23072 15660 23100
rect 15151 23069 15163 23072
rect 15105 23063 15163 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15197 23035 15255 23041
rect 11388 23004 14780 23032
rect 15028 23004 15148 23032
rect 11388 22992 11394 23004
rect 9585 22967 9643 22973
rect 9585 22933 9597 22967
rect 9631 22964 9643 22967
rect 10042 22964 10048 22976
rect 9631 22936 10048 22964
rect 9631 22933 9643 22936
rect 9585 22927 9643 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 11238 22924 11244 22976
rect 11296 22924 11302 22976
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12676 22936 13001 22964
rect 12676 22924 12682 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 13357 22967 13415 22973
rect 13357 22933 13369 22967
rect 13403 22964 13415 22967
rect 14458 22964 14464 22976
rect 13403 22936 14464 22964
rect 13403 22933 13415 22936
rect 13357 22927 13415 22933
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 14752 22973 14780 23004
rect 14737 22967 14795 22973
rect 14737 22933 14749 22967
rect 14783 22933 14795 22967
rect 15120 22964 15148 23004
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 15856 23032 15884 23267
rect 17310 23264 17316 23276
rect 17368 23304 17374 23316
rect 17368 23276 22094 23304
rect 17368 23264 17374 23276
rect 18601 23239 18659 23245
rect 18601 23205 18613 23239
rect 18647 23236 18659 23239
rect 19426 23236 19432 23248
rect 18647 23208 19432 23236
rect 18647 23205 18659 23208
rect 18601 23199 18659 23205
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 22066 23236 22094 23276
rect 25498 23264 25504 23316
rect 25556 23304 25562 23316
rect 26050 23304 26056 23316
rect 25556 23276 26056 23304
rect 25556 23264 25562 23276
rect 26050 23264 26056 23276
rect 26108 23264 26114 23316
rect 26418 23236 26424 23248
rect 22066 23208 26424 23236
rect 26418 23196 26424 23208
rect 26476 23196 26482 23248
rect 18049 23171 18107 23177
rect 18049 23137 18061 23171
rect 18095 23168 18107 23171
rect 18414 23168 18420 23180
rect 18095 23140 18420 23168
rect 18095 23137 18107 23140
rect 18049 23131 18107 23137
rect 18414 23128 18420 23140
rect 18472 23128 18478 23180
rect 18969 23171 19027 23177
rect 18969 23137 18981 23171
rect 19015 23168 19027 23171
rect 19058 23168 19064 23180
rect 19015 23140 19064 23168
rect 19015 23137 19027 23140
rect 18969 23131 19027 23137
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 20070 23128 20076 23180
rect 20128 23128 20134 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 20901 23171 20959 23177
rect 20901 23168 20913 23171
rect 20864 23140 20913 23168
rect 20864 23128 20870 23140
rect 20901 23137 20913 23140
rect 20947 23137 20959 23171
rect 20901 23131 20959 23137
rect 23385 23171 23443 23177
rect 23385 23137 23397 23171
rect 23431 23168 23443 23171
rect 24854 23168 24860 23180
rect 23431 23140 24860 23168
rect 23431 23137 23443 23140
rect 23385 23131 23443 23137
rect 24854 23128 24860 23140
rect 24912 23128 24918 23180
rect 24946 23128 24952 23180
rect 25004 23168 25010 23180
rect 25133 23171 25191 23177
rect 25133 23168 25145 23171
rect 25004 23140 25145 23168
rect 25004 23128 25010 23140
rect 25133 23137 25145 23140
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 18138 23060 18144 23112
rect 18196 23060 18202 23112
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 18598 23100 18604 23112
rect 18279 23072 18604 23100
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 18598 23060 18604 23072
rect 18656 23060 18662 23112
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20254 23100 20260 23112
rect 19935 23072 20260 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20254 23060 20260 23072
rect 20312 23060 20318 23112
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24026 23060 24032 23112
rect 24084 23100 24090 23112
rect 25041 23103 25099 23109
rect 25041 23100 25053 23103
rect 24084 23072 25053 23100
rect 24084 23060 24090 23072
rect 25041 23069 25053 23072
rect 25087 23069 25099 23103
rect 25041 23063 25099 23069
rect 15243 23004 15884 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 17862 22964 17868 22976
rect 15120 22936 17868 22964
rect 14737 22927 14795 22933
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 18156 22964 18184 23060
rect 18506 22992 18512 23044
rect 18564 23032 18570 23044
rect 22002 23032 22008 23044
rect 18564 23004 19564 23032
rect 18564 22992 18570 23004
rect 18690 22964 18696 22976
rect 18156 22936 18696 22964
rect 18690 22924 18696 22936
rect 18748 22924 18754 22976
rect 19536 22973 19564 23004
rect 19996 23004 22008 23032
rect 19996 22973 20024 23004
rect 22002 22992 22008 23004
rect 22060 22992 22066 23044
rect 24949 23035 25007 23041
rect 24949 23001 24961 23035
rect 24995 23032 25007 23035
rect 25130 23032 25136 23044
rect 24995 23004 25136 23032
rect 24995 23001 25007 23004
rect 24949 22995 25007 23001
rect 25130 22992 25136 23004
rect 25188 22992 25194 23044
rect 19521 22967 19579 22973
rect 19521 22933 19533 22967
rect 19567 22933 19579 22967
rect 19521 22927 19579 22933
rect 19981 22967 20039 22973
rect 19981 22933 19993 22967
rect 20027 22933 20039 22967
rect 19981 22927 20039 22933
rect 21821 22967 21879 22973
rect 21821 22933 21833 22967
rect 21867 22964 21879 22967
rect 22094 22964 22100 22976
rect 21867 22936 22100 22964
rect 21867 22933 21879 22936
rect 21821 22927 21879 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 24026 22924 24032 22976
rect 24084 22964 24090 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 24084 22936 24593 22964
rect 24084 22924 24090 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 7558 22720 7564 22772
rect 7616 22760 7622 22772
rect 8113 22763 8171 22769
rect 8113 22760 8125 22763
rect 7616 22732 8125 22760
rect 7616 22720 7622 22732
rect 8113 22729 8125 22732
rect 8159 22760 8171 22763
rect 8294 22760 8300 22772
rect 8159 22732 8300 22760
rect 8159 22729 8171 22732
rect 8113 22723 8171 22729
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 12802 22760 12808 22772
rect 12636 22732 12808 22760
rect 9582 22652 9588 22704
rect 9640 22652 9646 22704
rect 9674 22652 9680 22704
rect 9732 22692 9738 22704
rect 12636 22701 12664 22732
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 13004 22732 14412 22760
rect 12621 22695 12679 22701
rect 9732 22664 9904 22692
rect 9732 22652 9738 22664
rect 8294 22584 8300 22636
rect 8352 22624 8358 22636
rect 9876 22633 9904 22664
rect 12621 22661 12633 22695
rect 12667 22661 12679 22695
rect 12621 22655 12679 22661
rect 12710 22652 12716 22704
rect 12768 22692 12774 22704
rect 13004 22692 13032 22732
rect 14384 22692 14412 22732
rect 14458 22720 14464 22772
rect 14516 22760 14522 22772
rect 14826 22760 14832 22772
rect 14516 22732 14832 22760
rect 14516 22720 14522 22732
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 17037 22763 17095 22769
rect 17037 22729 17049 22763
rect 17083 22729 17095 22763
rect 17037 22723 17095 22729
rect 14553 22695 14611 22701
rect 14553 22692 14565 22695
rect 12768 22664 13110 22692
rect 14384 22664 14565 22692
rect 12768 22652 12774 22664
rect 14553 22661 14565 22664
rect 14599 22661 14611 22695
rect 17052 22692 17080 22723
rect 18598 22720 18604 22772
rect 18656 22760 18662 22772
rect 18693 22763 18751 22769
rect 18693 22760 18705 22763
rect 18656 22732 18705 22760
rect 18656 22720 18662 22732
rect 18693 22729 18705 22732
rect 18739 22729 18751 22763
rect 18693 22723 18751 22729
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19668 22732 19717 22760
rect 19668 22720 19674 22732
rect 19705 22729 19717 22732
rect 19751 22729 19763 22763
rect 19705 22723 19763 22729
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 24670 22760 24676 22772
rect 21223 22732 24676 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 21634 22692 21640 22704
rect 17052 22664 21640 22692
rect 14553 22655 14611 22661
rect 21634 22652 21640 22664
rect 21692 22652 21698 22704
rect 9861 22627 9919 22633
rect 8352 22610 8510 22624
rect 8352 22596 8524 22610
rect 8352 22584 8358 22596
rect 8496 22556 8524 22596
rect 9861 22593 9873 22627
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 13906 22584 13912 22636
rect 13964 22624 13970 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 13964 22596 16865 22624
rect 13964 22584 13970 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 18690 22584 18696 22636
rect 18748 22624 18754 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18748 22596 18889 22624
rect 18748 22584 18754 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 20438 22584 20444 22636
rect 20496 22624 20502 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20496 22596 21097 22624
rect 20496 22584 20502 22596
rect 21085 22593 21097 22596
rect 21131 22624 21143 22627
rect 21450 22624 21456 22636
rect 21131 22596 21456 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 21450 22584 21456 22596
rect 21508 22584 21514 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 23934 22584 23940 22636
rect 23992 22584 23998 22636
rect 10137 22559 10195 22565
rect 10137 22556 10149 22559
rect 8496 22528 10149 22556
rect 10137 22525 10149 22528
rect 10183 22525 10195 22559
rect 10137 22519 10195 22525
rect 19702 22516 19708 22568
rect 19760 22556 19766 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 19760 22528 21281 22556
rect 19760 22516 19766 22528
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 22830 22516 22836 22568
rect 22888 22516 22894 22568
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 9784 22460 12434 22488
rect 9398 22380 9404 22432
rect 9456 22420 9462 22432
rect 9784 22420 9812 22460
rect 9456 22392 9812 22420
rect 12406 22420 12434 22460
rect 18598 22448 18604 22500
rect 18656 22488 18662 22500
rect 20806 22488 20812 22500
rect 18656 22460 20812 22488
rect 18656 22448 18662 22460
rect 20806 22448 20812 22460
rect 20864 22448 20870 22500
rect 12986 22420 12992 22432
rect 12406 22392 12992 22420
rect 9456 22380 9462 22392
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 20438 22380 20444 22432
rect 20496 22380 20502 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 15930 22216 15936 22228
rect 9824 22188 15936 22216
rect 9824 22176 9830 22188
rect 15930 22176 15936 22188
rect 15988 22176 15994 22228
rect 18690 22176 18696 22228
rect 18748 22216 18754 22228
rect 21082 22216 21088 22228
rect 18748 22188 21088 22216
rect 18748 22176 18754 22188
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 23753 22219 23811 22225
rect 23753 22185 23765 22219
rect 23799 22216 23811 22219
rect 23842 22216 23848 22228
rect 23799 22188 23848 22216
rect 23799 22185 23811 22188
rect 23753 22179 23811 22185
rect 23842 22176 23848 22188
rect 23900 22176 23906 22228
rect 25406 22216 25412 22228
rect 25148 22188 25412 22216
rect 6914 22108 6920 22160
rect 6972 22148 6978 22160
rect 7834 22148 7840 22160
rect 6972 22120 7840 22148
rect 6972 22108 6978 22120
rect 7834 22108 7840 22120
rect 7892 22148 7898 22160
rect 9674 22148 9680 22160
rect 7892 22120 9680 22148
rect 7892 22108 7898 22120
rect 9674 22108 9680 22120
rect 9732 22108 9738 22160
rect 11054 22148 11060 22160
rect 10888 22120 11060 22148
rect 10888 22089 10916 22120
rect 11054 22108 11060 22120
rect 11112 22108 11118 22160
rect 11146 22108 11152 22160
rect 11204 22148 11210 22160
rect 12526 22148 12532 22160
rect 11204 22120 12112 22148
rect 11204 22108 11210 22120
rect 12084 22089 12112 22120
rect 12268 22120 12532 22148
rect 12268 22089 12296 22120
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 15746 22148 15752 22160
rect 15120 22120 15752 22148
rect 10873 22083 10931 22089
rect 10873 22049 10885 22083
rect 10919 22049 10931 22083
rect 10873 22043 10931 22049
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22049 12127 22083
rect 12069 22043 12127 22049
rect 12253 22083 12311 22089
rect 12253 22049 12265 22083
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 14090 22040 14096 22092
rect 14148 22080 14154 22092
rect 14550 22080 14556 22092
rect 14148 22052 14556 22080
rect 14148 22040 14154 22052
rect 14550 22040 14556 22052
rect 14608 22080 14614 22092
rect 15120 22089 15148 22120
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 17862 22108 17868 22160
rect 17920 22108 17926 22160
rect 14921 22083 14979 22089
rect 14921 22080 14933 22083
rect 14608 22052 14933 22080
rect 14608 22040 14614 22052
rect 14921 22049 14933 22052
rect 14967 22049 14979 22083
rect 14921 22043 14979 22049
rect 15105 22083 15163 22089
rect 15105 22049 15117 22083
rect 15151 22080 15163 22083
rect 16117 22083 16175 22089
rect 15151 22052 15185 22080
rect 15151 22049 15163 22052
rect 15105 22043 15163 22049
rect 16117 22049 16129 22083
rect 16163 22080 16175 22083
rect 16942 22080 16948 22092
rect 16163 22052 16948 22080
rect 16163 22049 16175 22052
rect 16117 22043 16175 22049
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 17880 22080 17908 22108
rect 19058 22080 19064 22092
rect 17880 22052 19064 22080
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 19889 22083 19947 22089
rect 19889 22049 19901 22083
rect 19935 22080 19947 22083
rect 20622 22080 20628 22092
rect 19935 22052 20628 22080
rect 19935 22049 19947 22052
rect 19889 22043 19947 22049
rect 20622 22040 20628 22052
rect 20680 22040 20686 22092
rect 25148 22089 25176 22188
rect 25406 22176 25412 22188
rect 25464 22176 25470 22228
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22080 21143 22083
rect 25133 22083 25191 22089
rect 21131 22052 24992 22080
rect 21131 22049 21143 22052
rect 21085 22043 21143 22049
rect 21542 21972 21548 22024
rect 21600 22012 21606 22024
rect 21600 21984 21942 22012
rect 21600 21972 21606 21984
rect 23290 21972 23296 22024
rect 23348 21972 23354 22024
rect 24964 22021 24992 22052
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 22012 25099 22015
rect 25222 22012 25228 22024
rect 25087 21984 25228 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 11146 21904 11152 21956
rect 11204 21944 11210 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 11204 21916 12357 21944
rect 11204 21904 11210 21916
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12345 21907 12403 21913
rect 15930 21904 15936 21956
rect 15988 21944 15994 21956
rect 16393 21947 16451 21953
rect 16393 21944 16405 21947
rect 15988 21916 16405 21944
rect 15988 21904 15994 21916
rect 16393 21913 16405 21916
rect 16439 21944 16451 21947
rect 16482 21944 16488 21956
rect 16439 21916 16488 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 16482 21904 16488 21916
rect 16540 21904 16546 21956
rect 18233 21947 18291 21953
rect 18233 21944 18245 21947
rect 17618 21916 18245 21944
rect 8294 21836 8300 21888
rect 8352 21876 8358 21888
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8352 21848 8953 21876
rect 8352 21836 8358 21848
rect 8941 21845 8953 21848
rect 8987 21845 8999 21879
rect 8941 21839 8999 21845
rect 10413 21879 10471 21885
rect 10413 21845 10425 21879
rect 10459 21876 10471 21879
rect 10594 21876 10600 21888
rect 10459 21848 10600 21876
rect 10459 21845 10471 21848
rect 10413 21839 10471 21845
rect 10594 21836 10600 21848
rect 10652 21876 10658 21888
rect 10965 21879 11023 21885
rect 10965 21876 10977 21879
rect 10652 21848 10977 21876
rect 10652 21836 10658 21848
rect 10965 21845 10977 21848
rect 11011 21845 11023 21879
rect 10965 21839 11023 21845
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 11422 21836 11428 21888
rect 11480 21836 11486 21888
rect 12713 21879 12771 21885
rect 12713 21845 12725 21879
rect 12759 21876 12771 21879
rect 13906 21876 13912 21888
rect 12759 21848 13912 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 13906 21836 13912 21848
rect 13964 21836 13970 21888
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 15197 21879 15255 21885
rect 15197 21876 15209 21879
rect 14056 21848 15209 21876
rect 14056 21836 14062 21848
rect 15197 21845 15209 21848
rect 15243 21845 15255 21879
rect 15197 21839 15255 21845
rect 15565 21879 15623 21885
rect 15565 21845 15577 21879
rect 15611 21876 15623 21879
rect 15838 21876 15844 21888
rect 15611 21848 15844 21876
rect 15611 21845 15623 21848
rect 15565 21839 15623 21845
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 17402 21836 17408 21888
rect 17460 21876 17466 21888
rect 17696 21876 17724 21916
rect 18233 21913 18245 21916
rect 18279 21913 18291 21947
rect 18233 21907 18291 21913
rect 23014 21904 23020 21956
rect 23072 21904 23078 21956
rect 17460 21848 17724 21876
rect 17460 21836 17466 21848
rect 17862 21836 17868 21888
rect 17920 21836 17926 21888
rect 19610 21836 19616 21888
rect 19668 21876 19674 21888
rect 19978 21876 19984 21888
rect 19668 21848 19984 21876
rect 19668 21836 19674 21848
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 20070 21836 20076 21888
rect 20128 21836 20134 21888
rect 20346 21836 20352 21888
rect 20404 21876 20410 21888
rect 20441 21879 20499 21885
rect 20441 21876 20453 21879
rect 20404 21848 20453 21876
rect 20404 21836 20410 21848
rect 20441 21845 20453 21848
rect 20487 21845 20499 21879
rect 20441 21839 20499 21845
rect 20898 21836 20904 21888
rect 20956 21876 20962 21888
rect 21545 21879 21603 21885
rect 21545 21876 21557 21879
rect 20956 21848 21557 21876
rect 20956 21836 20962 21848
rect 21545 21845 21557 21848
rect 21591 21845 21603 21879
rect 21545 21839 21603 21845
rect 22002 21836 22008 21888
rect 22060 21876 22066 21888
rect 23952 21876 23980 21975
rect 25222 21972 25228 21984
rect 25280 21972 25286 22024
rect 22060 21848 23980 21876
rect 22060 21836 22066 21848
rect 24394 21836 24400 21888
rect 24452 21876 24458 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 24452 21848 24593 21876
rect 24452 21836 24458 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 8662 21632 8668 21684
rect 8720 21632 8726 21684
rect 9950 21632 9956 21684
rect 10008 21632 10014 21684
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11112 21644 11713 21672
rect 11112 21632 11118 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 12710 21632 12716 21684
rect 12768 21672 12774 21684
rect 15102 21672 15108 21684
rect 12768 21644 15108 21672
rect 12768 21632 12774 21644
rect 10873 21607 10931 21613
rect 10873 21573 10885 21607
rect 10919 21604 10931 21607
rect 12158 21604 12164 21616
rect 10919 21576 12164 21604
rect 10919 21573 10931 21576
rect 10873 21567 10931 21573
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 14200 21604 14228 21644
rect 15102 21632 15108 21644
rect 15160 21632 15166 21684
rect 18690 21632 18696 21684
rect 18748 21672 18754 21684
rect 19797 21675 19855 21681
rect 19797 21672 19809 21675
rect 18748 21644 19809 21672
rect 18748 21632 18754 21644
rect 19797 21641 19809 21644
rect 19843 21641 19855 21675
rect 19797 21635 19855 21641
rect 20070 21632 20076 21684
rect 20128 21672 20134 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20128 21644 21189 21672
rect 20128 21632 20134 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22554 21672 22560 21684
rect 22511 21644 22560 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 23348 21644 25084 21672
rect 23348 21632 23354 21644
rect 14122 21576 14228 21604
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 15749 21607 15807 21613
rect 14332 21576 14872 21604
rect 14332 21564 14338 21576
rect 8294 21496 8300 21548
rect 8352 21496 8358 21548
rect 9214 21496 9220 21548
rect 9272 21536 9278 21548
rect 9493 21539 9551 21545
rect 9493 21536 9505 21539
rect 9272 21508 9505 21536
rect 9272 21496 9278 21508
rect 9493 21505 9505 21508
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9950 21536 9956 21548
rect 9631 21508 9956 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 11606 21536 11612 21548
rect 10827 21508 11612 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 14844 21545 14872 21576
rect 15749 21573 15761 21607
rect 15795 21604 15807 21607
rect 18782 21604 18788 21616
rect 15795 21576 18788 21604
rect 15795 21573 15807 21576
rect 15749 21567 15807 21573
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 21361 21607 21419 21613
rect 21361 21604 21373 21607
rect 20036 21576 21373 21604
rect 20036 21564 20042 21576
rect 21361 21573 21373 21576
rect 21407 21573 21419 21607
rect 21361 21567 21419 21573
rect 21542 21564 21548 21616
rect 21600 21604 21606 21616
rect 21600 21590 23598 21604
rect 21600 21576 23612 21590
rect 21600 21564 21606 21576
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 15896 21508 18705 21536
rect 15896 21496 15902 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 19935 21508 20729 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20717 21505 20729 21508
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22244 21508 22385 21536
rect 22244 21496 22250 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 23584 21480 23612 21576
rect 25056 21545 25084 21644
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21505 25099 21539
rect 25041 21499 25099 21505
rect 6914 21428 6920 21480
rect 6972 21428 6978 21480
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 7742 21468 7748 21480
rect 7239 21440 7748 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 7742 21428 7748 21440
rect 7800 21428 7806 21480
rect 9306 21428 9312 21480
rect 9364 21428 9370 21480
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 19702 21428 19708 21480
rect 19760 21428 19766 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 23474 21468 23480 21480
rect 22695 21440 23480 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 23566 21428 23572 21480
rect 23624 21428 23630 21480
rect 24394 21468 24400 21480
rect 23768 21440 24400 21468
rect 15562 21360 15568 21412
rect 15620 21360 15626 21412
rect 18877 21403 18935 21409
rect 18877 21369 18889 21403
rect 18923 21400 18935 21403
rect 21634 21400 21640 21412
rect 18923 21372 21640 21400
rect 18923 21369 18935 21372
rect 18877 21363 18935 21369
rect 21634 21360 21640 21372
rect 21692 21360 21698 21412
rect 22830 21360 22836 21412
rect 22888 21400 22894 21412
rect 23768 21400 23796 21440
rect 24394 21428 24400 21440
rect 24452 21428 24458 21480
rect 24765 21471 24823 21477
rect 24765 21437 24777 21471
rect 24811 21468 24823 21471
rect 25314 21468 25320 21480
rect 24811 21440 25320 21468
rect 24811 21437 24823 21440
rect 24765 21431 24823 21437
rect 22888 21372 23796 21400
rect 22888 21360 22894 21372
rect 24964 21344 24992 21440
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 13081 21335 13139 21341
rect 13081 21332 13093 21335
rect 12768 21304 13093 21332
rect 12768 21292 12774 21304
rect 13081 21301 13093 21304
rect 13127 21332 13139 21335
rect 13538 21332 13544 21344
rect 13127 21304 13544 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 15102 21292 15108 21344
rect 15160 21292 15166 21344
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 19153 21335 19211 21341
rect 19153 21332 19165 21335
rect 18840 21304 19165 21332
rect 18840 21292 18846 21304
rect 19153 21301 19165 21304
rect 19199 21301 19211 21335
rect 19153 21295 19211 21301
rect 20257 21335 20315 21341
rect 20257 21301 20269 21335
rect 20303 21332 20315 21335
rect 20438 21332 20444 21344
rect 20303 21304 20444 21332
rect 20303 21301 20315 21304
rect 20257 21295 20315 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21542 21292 21548 21344
rect 21600 21292 21606 21344
rect 22002 21292 22008 21344
rect 22060 21292 22066 21344
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23290 21332 23296 21344
rect 23072 21304 23296 21332
rect 23072 21292 23078 21304
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 24946 21292 24952 21344
rect 25004 21292 25010 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 21082 21088 21088 21140
rect 21140 21128 21146 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 21140 21100 21465 21128
rect 21140 21088 21146 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 21453 21091 21511 21097
rect 20993 21063 21051 21069
rect 12084 21032 12940 21060
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 10689 20995 10747 21001
rect 10689 20992 10701 20995
rect 9732 20964 10701 20992
rect 9732 20952 9738 20964
rect 10689 20961 10701 20964
rect 10735 20961 10747 20995
rect 10689 20955 10747 20961
rect 12084 20936 12112 21032
rect 9950 20884 9956 20936
rect 10008 20884 10014 20936
rect 12066 20884 12072 20936
rect 12124 20884 12130 20936
rect 10962 20816 10968 20868
rect 11020 20816 11026 20868
rect 12802 20856 12808 20868
rect 12544 20828 12808 20856
rect 12544 20800 12572 20828
rect 12802 20816 12808 20828
rect 12860 20816 12866 20868
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9214 20788 9220 20800
rect 9171 20760 9220 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9214 20748 9220 20760
rect 9272 20748 9278 20800
rect 12437 20791 12495 20797
rect 12437 20757 12449 20791
rect 12483 20788 12495 20791
rect 12526 20788 12532 20800
rect 12483 20760 12532 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 12713 20791 12771 20797
rect 12713 20757 12725 20791
rect 12759 20788 12771 20791
rect 12912 20788 12940 21032
rect 16868 21032 20852 21060
rect 15194 20952 15200 21004
rect 15252 20992 15258 21004
rect 16868 20992 16896 21032
rect 15252 20964 16896 20992
rect 15252 20952 15258 20964
rect 16942 20952 16948 21004
rect 17000 20952 17006 21004
rect 19610 20952 19616 21004
rect 19668 20952 19674 21004
rect 17218 20884 17224 20936
rect 17276 20924 17282 20936
rect 17770 20924 17776 20936
rect 17276 20896 17776 20924
rect 17276 20884 17282 20896
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 20824 20933 20852 21032
rect 20993 21029 21005 21063
rect 21039 21060 21051 21063
rect 21039 21032 22094 21060
rect 21039 21029 21051 21032
rect 20993 21023 21051 21029
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19300 20896 19809 20924
rect 19300 20884 19306 20896
rect 19797 20893 19809 20896
rect 19843 20924 19855 20927
rect 20441 20927 20499 20933
rect 20441 20924 20453 20927
rect 19843 20896 20453 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 20441 20893 20453 20896
rect 20487 20893 20499 20927
rect 20441 20887 20499 20893
rect 20809 20927 20867 20933
rect 20809 20893 20821 20927
rect 20855 20893 20867 20927
rect 22066 20924 22094 21032
rect 22186 20952 22192 21004
rect 22244 20952 22250 21004
rect 24670 20952 24676 21004
rect 24728 20952 24734 21004
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25406 20992 25412 21004
rect 25004 20964 25412 20992
rect 25004 20952 25010 20964
rect 25406 20952 25412 20964
rect 25464 20952 25470 21004
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22066 20896 22661 20924
rect 20809 20887 20867 20893
rect 22649 20893 22661 20896
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20924 23903 20927
rect 24854 20924 24860 20936
rect 23891 20896 24860 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 25038 20884 25044 20936
rect 25096 20884 25102 20936
rect 14660 20828 15502 20856
rect 14660 20800 14688 20828
rect 16574 20816 16580 20868
rect 16632 20856 16638 20868
rect 16669 20859 16727 20865
rect 16669 20856 16681 20859
rect 16632 20828 16681 20856
rect 16632 20816 16638 20828
rect 16669 20825 16681 20828
rect 16715 20825 16727 20859
rect 16669 20819 16727 20825
rect 19058 20816 19064 20868
rect 19116 20856 19122 20868
rect 19705 20859 19763 20865
rect 19705 20856 19717 20859
rect 19116 20828 19717 20856
rect 19116 20816 19122 20828
rect 19705 20825 19717 20828
rect 19751 20856 19763 20859
rect 21269 20859 21327 20865
rect 21269 20856 21281 20859
rect 19751 20828 21281 20856
rect 19751 20825 19763 20828
rect 19705 20819 19763 20825
rect 21269 20825 21281 20828
rect 21315 20825 21327 20859
rect 25056 20856 25084 20884
rect 21269 20819 21327 20825
rect 24872 20828 25084 20856
rect 14642 20788 14648 20800
rect 12759 20760 14648 20788
rect 12759 20757 12771 20760
rect 12713 20751 12771 20757
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 15197 20791 15255 20797
rect 15197 20757 15209 20791
rect 15243 20788 15255 20791
rect 15838 20788 15844 20800
rect 15243 20760 15844 20788
rect 15243 20757 15255 20760
rect 15197 20751 15255 20757
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17402 20788 17408 20800
rect 17276 20760 17408 20788
rect 17276 20748 17282 20760
rect 17402 20748 17408 20760
rect 17460 20788 17466 20800
rect 18693 20791 18751 20797
rect 18693 20788 18705 20791
rect 17460 20760 18705 20788
rect 17460 20748 17466 20760
rect 18693 20757 18705 20760
rect 18739 20757 18751 20791
rect 18693 20751 18751 20757
rect 19886 20748 19892 20800
rect 19944 20788 19950 20800
rect 24872 20797 24900 20828
rect 20165 20791 20223 20797
rect 20165 20788 20177 20791
rect 19944 20760 20177 20788
rect 19944 20748 19950 20760
rect 20165 20757 20177 20760
rect 20211 20757 20223 20791
rect 20165 20751 20223 20757
rect 24857 20791 24915 20797
rect 24857 20757 24869 20791
rect 24903 20757 24915 20791
rect 24857 20751 24915 20757
rect 24946 20748 24952 20800
rect 25004 20748 25010 20800
rect 25038 20748 25044 20800
rect 25096 20788 25102 20800
rect 25317 20791 25375 20797
rect 25317 20788 25329 20791
rect 25096 20760 25329 20788
rect 25096 20748 25102 20760
rect 25317 20757 25329 20760
rect 25363 20757 25375 20791
rect 25317 20751 25375 20757
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 10045 20587 10103 20593
rect 10045 20584 10057 20587
rect 8404 20556 10057 20584
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 8404 20516 8432 20556
rect 10045 20553 10057 20556
rect 10091 20553 10103 20587
rect 10045 20547 10103 20553
rect 10410 20544 10416 20596
rect 10468 20544 10474 20596
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 11330 20584 11336 20596
rect 10827 20556 11336 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 15378 20584 15384 20596
rect 15335 20556 15384 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 16758 20544 16764 20596
rect 16816 20584 16822 20596
rect 18414 20584 18420 20596
rect 16816 20556 18420 20584
rect 16816 20544 16822 20556
rect 18414 20544 18420 20556
rect 18472 20544 18478 20596
rect 21726 20584 21732 20596
rect 20456 20556 21732 20584
rect 14642 20516 14648 20528
rect 8352 20488 8510 20516
rect 14214 20488 14648 20516
rect 8352 20476 8358 20488
rect 14642 20476 14648 20488
rect 14700 20516 14706 20528
rect 15102 20516 15108 20528
rect 14700 20488 15108 20516
rect 14700 20476 14706 20488
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 20162 20516 20168 20528
rect 19260 20488 20168 20516
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 6914 20448 6920 20460
rect 6604 20420 6920 20448
rect 6604 20408 6610 20420
rect 6914 20408 6920 20420
rect 6972 20448 6978 20460
rect 7745 20451 7803 20457
rect 7745 20448 7757 20451
rect 6972 20420 7757 20448
rect 6972 20408 6978 20420
rect 7745 20417 7757 20420
rect 7791 20417 7803 20451
rect 7745 20411 7803 20417
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 12492 20420 12725 20448
rect 12492 20408 12498 20420
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20448 18659 20451
rect 19150 20448 19156 20460
rect 18647 20420 19156 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 19260 20457 19288 20488
rect 20162 20476 20168 20488
rect 20220 20476 20226 20528
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20456 20448 20484 20556
rect 21726 20544 21732 20556
rect 21784 20544 21790 20596
rect 23293 20587 23351 20593
rect 23293 20553 23305 20587
rect 23339 20584 23351 20587
rect 23566 20584 23572 20596
rect 23339 20556 23572 20584
rect 23339 20553 23351 20556
rect 23293 20547 23351 20553
rect 23566 20544 23572 20556
rect 23624 20584 23630 20596
rect 23842 20584 23848 20596
rect 23624 20556 23848 20584
rect 23624 20544 23630 20556
rect 23842 20544 23848 20556
rect 23900 20544 23906 20596
rect 25314 20544 25320 20596
rect 25372 20544 25378 20596
rect 20806 20476 20812 20528
rect 20864 20516 20870 20528
rect 21453 20519 21511 20525
rect 21453 20516 21465 20519
rect 20864 20488 21465 20516
rect 20864 20476 20870 20488
rect 21453 20485 21465 20488
rect 21499 20485 21511 20519
rect 21453 20479 21511 20485
rect 21634 20476 21640 20528
rect 21692 20516 21698 20528
rect 23860 20516 23888 20544
rect 21692 20488 22784 20516
rect 23860 20488 24334 20516
rect 21692 20476 21698 20488
rect 22756 20457 22784 20488
rect 19935 20420 20484 20448
rect 22005 20451 22063 20457
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22741 20451 22799 20457
rect 22741 20417 22753 20451
rect 22787 20417 22799 20451
rect 22741 20411 22799 20417
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8662 20380 8668 20392
rect 8067 20352 8668 20380
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8662 20340 8668 20352
rect 8720 20340 8726 20392
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 10134 20380 10140 20392
rect 9815 20352 10140 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 10410 20340 10416 20392
rect 10468 20380 10474 20392
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10468 20352 10885 20380
rect 10468 20340 10474 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 10965 20343 11023 20349
rect 12728 20352 13001 20380
rect 10778 20272 10784 20324
rect 10836 20312 10842 20324
rect 10980 20312 11008 20343
rect 12728 20324 12756 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 15105 20383 15163 20389
rect 15105 20380 15117 20383
rect 12989 20343 13047 20349
rect 14476 20352 15117 20380
rect 10836 20284 11008 20312
rect 10836 20272 10842 20284
rect 12710 20272 12716 20324
rect 12768 20272 12774 20324
rect 14476 20256 14504 20352
rect 15105 20349 15117 20352
rect 15151 20349 15163 20383
rect 15105 20343 15163 20349
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 18325 20383 18383 20389
rect 18325 20380 18337 20383
rect 17920 20352 18337 20380
rect 17920 20340 17926 20352
rect 18325 20349 18337 20352
rect 18371 20349 18383 20383
rect 18325 20343 18383 20349
rect 20530 20340 20536 20392
rect 20588 20340 20594 20392
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 21082 20380 21088 20392
rect 20763 20352 21088 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 21082 20340 21088 20352
rect 21140 20340 21146 20392
rect 22020 20312 22048 20411
rect 23566 20340 23572 20392
rect 23624 20340 23630 20392
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 25130 20380 25136 20392
rect 23891 20352 25136 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 18524 20284 22048 20312
rect 22189 20315 22247 20321
rect 14458 20204 14464 20256
rect 14516 20204 14522 20256
rect 15746 20204 15752 20256
rect 15804 20204 15810 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 16853 20247 16911 20253
rect 16853 20244 16865 20247
rect 16816 20216 16865 20244
rect 16816 20204 16822 20216
rect 16853 20213 16865 20216
rect 16899 20213 16911 20247
rect 16853 20207 16911 20213
rect 17034 20204 17040 20256
rect 17092 20244 17098 20256
rect 18524 20244 18552 20284
rect 22189 20281 22201 20315
rect 22235 20312 22247 20315
rect 23474 20312 23480 20324
rect 22235 20284 23480 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 17092 20216 18552 20244
rect 17092 20204 17098 20216
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 19702 20204 19708 20256
rect 19760 20204 19766 20256
rect 21177 20247 21235 20253
rect 21177 20213 21189 20247
rect 21223 20244 21235 20247
rect 21726 20244 21732 20256
rect 21223 20216 21732 20244
rect 21223 20213 21235 20216
rect 21177 20207 21235 20213
rect 21726 20204 21732 20216
rect 21784 20204 21790 20256
rect 22738 20204 22744 20256
rect 22796 20244 22802 20256
rect 22925 20247 22983 20253
rect 22925 20244 22937 20247
rect 22796 20216 22937 20244
rect 22796 20204 22802 20216
rect 22925 20213 22937 20216
rect 22971 20213 22983 20247
rect 22925 20207 22983 20213
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 10873 20043 10931 20049
rect 10873 20009 10885 20043
rect 10919 20040 10931 20043
rect 10962 20040 10968 20052
rect 10919 20012 10968 20040
rect 10919 20009 10931 20012
rect 10873 20003 10931 20009
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 12069 20043 12127 20049
rect 12069 20009 12081 20043
rect 12115 20040 12127 20043
rect 13354 20040 13360 20052
rect 12115 20012 13360 20040
rect 12115 20009 12127 20012
rect 12069 20003 12127 20009
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 15102 20000 15108 20052
rect 15160 20040 15166 20052
rect 16025 20043 16083 20049
rect 15160 20012 15976 20040
rect 15160 20000 15166 20012
rect 15948 19972 15976 20012
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16574 20040 16580 20052
rect 16071 20012 16580 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 16669 20043 16727 20049
rect 16669 20009 16681 20043
rect 16715 20040 16727 20043
rect 17034 20040 17040 20052
rect 16715 20012 17040 20040
rect 16715 20009 16727 20012
rect 16669 20003 16727 20009
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 18233 20043 18291 20049
rect 18233 20009 18245 20043
rect 18279 20040 18291 20043
rect 21174 20040 21180 20052
rect 18279 20012 21180 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 21174 20000 21180 20012
rect 21232 20000 21238 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 23845 20043 23903 20049
rect 23845 20040 23857 20043
rect 23716 20012 23857 20040
rect 23716 20000 23722 20012
rect 23845 20009 23857 20012
rect 23891 20040 23903 20043
rect 24670 20040 24676 20052
rect 23891 20012 24676 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 16945 19975 17003 19981
rect 16945 19972 16957 19975
rect 15948 19944 16957 19972
rect 16945 19941 16957 19944
rect 16991 19972 17003 19975
rect 17218 19972 17224 19984
rect 16991 19944 17224 19972
rect 16991 19941 17003 19944
rect 16945 19935 17003 19941
rect 17218 19932 17224 19944
rect 17276 19932 17282 19984
rect 9398 19864 9404 19916
rect 9456 19864 9462 19916
rect 11514 19864 11520 19916
rect 11572 19864 11578 19916
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 13354 19904 13360 19916
rect 12492 19876 13360 19904
rect 12492 19864 12498 19876
rect 13354 19864 13360 19876
rect 13412 19904 13418 19916
rect 14274 19904 14280 19916
rect 13412 19876 14280 19904
rect 13412 19864 13418 19876
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 14550 19864 14556 19916
rect 14608 19904 14614 19916
rect 17681 19907 17739 19913
rect 14608 19876 16528 19904
rect 14608 19864 14614 19876
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 16500 19845 16528 19876
rect 17681 19873 17693 19907
rect 17727 19904 17739 19907
rect 17862 19904 17868 19916
rect 17727 19876 17868 19904
rect 17727 19873 17739 19876
rect 17681 19867 17739 19873
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 20254 19904 20260 19916
rect 19935 19876 20260 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 20254 19864 20260 19876
rect 20312 19904 20318 19916
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 20312 19876 22109 19904
rect 20312 19864 20318 19876
rect 22097 19873 22109 19876
rect 22143 19873 22155 19907
rect 22097 19867 22155 19873
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19836 17831 19839
rect 18322 19836 18328 19848
rect 17819 19808 18328 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19836 18935 19839
rect 19518 19836 19524 19848
rect 18923 19808 19524 19836
rect 18923 19805 18935 19808
rect 18877 19799 18935 19805
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 14553 19771 14611 19777
rect 8404 19740 9890 19768
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 8404 19709 8432 19740
rect 9600 19712 9628 19740
rect 14553 19737 14565 19771
rect 14599 19768 14611 19771
rect 14826 19768 14832 19780
rect 14599 19740 14832 19768
rect 14599 19737 14611 19740
rect 14553 19731 14611 19737
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 15102 19728 15108 19780
rect 15160 19728 15166 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 16592 19740 17877 19768
rect 8389 19703 8447 19709
rect 8389 19700 8401 19703
rect 8352 19672 8401 19700
rect 8352 19660 8358 19672
rect 8389 19669 8401 19672
rect 8435 19669 8447 19703
rect 8389 19663 8447 19669
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 11422 19660 11428 19712
rect 11480 19700 11486 19712
rect 11609 19703 11667 19709
rect 11609 19700 11621 19703
rect 11480 19672 11621 19700
rect 11480 19660 11486 19672
rect 11609 19669 11621 19672
rect 11655 19669 11667 19703
rect 11609 19663 11667 19669
rect 11698 19660 11704 19712
rect 11756 19660 11762 19712
rect 16482 19660 16488 19712
rect 16540 19700 16546 19712
rect 16592 19700 16620 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 17865 19731 17923 19737
rect 19794 19728 19800 19780
rect 19852 19768 19858 19780
rect 20162 19768 20168 19780
rect 19852 19740 20168 19768
rect 19852 19728 19858 19740
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 21542 19768 21548 19780
rect 21390 19740 21548 19768
rect 21542 19728 21548 19740
rect 21600 19728 21606 19780
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 22066 19740 22385 19768
rect 16540 19672 16620 19700
rect 16540 19660 16546 19672
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 22066 19700 22094 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 23842 19768 23848 19780
rect 23598 19740 23848 19768
rect 22373 19731 22431 19737
rect 23842 19728 23848 19740
rect 23900 19768 23906 19780
rect 24118 19768 24124 19780
rect 23900 19740 24124 19768
rect 23900 19728 23906 19740
rect 24118 19728 24124 19740
rect 24176 19768 24182 19780
rect 24397 19771 24455 19777
rect 24397 19768 24409 19771
rect 24176 19740 24409 19768
rect 24176 19728 24182 19740
rect 24397 19737 24409 19740
rect 24443 19768 24455 19771
rect 24581 19771 24639 19777
rect 24581 19768 24593 19771
rect 24443 19740 24593 19768
rect 24443 19737 24455 19740
rect 24397 19731 24455 19737
rect 24581 19737 24593 19740
rect 24627 19737 24639 19771
rect 24581 19731 24639 19737
rect 21692 19672 22094 19700
rect 24857 19703 24915 19709
rect 21692 19660 21698 19672
rect 24857 19669 24869 19703
rect 24903 19700 24915 19703
rect 24946 19700 24952 19712
rect 24903 19672 24952 19700
rect 24903 19669 24915 19672
rect 24857 19663 24915 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 9640 19468 10977 19496
rect 9640 19456 9646 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12529 19499 12587 19505
rect 12529 19496 12541 19499
rect 12492 19468 12541 19496
rect 12492 19456 12498 19468
rect 12529 19465 12541 19468
rect 12575 19465 12587 19499
rect 12529 19459 12587 19465
rect 15194 19456 15200 19508
rect 15252 19456 15258 19508
rect 17126 19456 17132 19508
rect 17184 19456 17190 19508
rect 17589 19499 17647 19505
rect 17589 19465 17601 19499
rect 17635 19496 17647 19499
rect 19242 19496 19248 19508
rect 17635 19468 19248 19496
rect 17635 19465 17647 19468
rect 17589 19459 17647 19465
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20438 19456 20444 19508
rect 20496 19456 20502 19508
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20714 19496 20720 19508
rect 20579 19468 20720 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 22189 19499 22247 19505
rect 22189 19465 22201 19499
rect 22235 19496 22247 19499
rect 22462 19496 22468 19508
rect 22235 19468 22468 19496
rect 22235 19465 22247 19468
rect 22189 19459 22247 19465
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 22649 19499 22707 19505
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 24026 19496 24032 19508
rect 22695 19468 24032 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 24026 19456 24032 19468
rect 24084 19456 24090 19508
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 8202 19428 8208 19440
rect 8050 19400 8208 19428
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 13906 19428 13912 19440
rect 13570 19400 13912 19428
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 14001 19431 14059 19437
rect 14001 19397 14013 19431
rect 14047 19428 14059 19431
rect 14458 19428 14464 19440
rect 14047 19400 14464 19428
rect 14047 19397 14059 19400
rect 14001 19391 14059 19397
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 15746 19388 15752 19440
rect 15804 19428 15810 19440
rect 22094 19428 22100 19440
rect 15804 19400 19012 19428
rect 15804 19388 15810 19400
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 9088 19332 9137 19360
rect 9088 19320 9094 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9950 19360 9956 19372
rect 9263 19332 9956 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 14274 19320 14280 19372
rect 14332 19320 14338 19372
rect 15010 19320 15016 19372
rect 15068 19320 15074 19372
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19360 16175 19363
rect 16390 19360 16396 19372
rect 16163 19332 16396 19360
rect 16163 19329 16175 19332
rect 16117 19323 16175 19329
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 18984 19369 19012 19400
rect 20640 19400 22100 19428
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17092 19332 17233 19360
rect 17092 19320 17098 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20640 19360 20668 19400
rect 22094 19388 22100 19400
rect 22152 19388 22158 19440
rect 23566 19428 23572 19440
rect 23400 19400 23572 19428
rect 23400 19369 23428 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 23658 19388 23664 19440
rect 23716 19388 23722 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 20588 19332 20668 19360
rect 21453 19363 21511 19369
rect 20588 19320 20594 19332
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 21499 19332 22569 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 6546 19252 6552 19304
rect 6604 19252 6610 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 6914 19292 6920 19304
rect 6871 19264 6920 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 6914 19252 6920 19264
rect 6972 19292 6978 19304
rect 7558 19292 7564 19304
rect 6972 19264 7564 19292
rect 6972 19252 6978 19264
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 8720 19264 9321 19292
rect 8720 19252 8726 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 9398 19252 9404 19304
rect 9456 19292 9462 19304
rect 9456 19264 16528 19292
rect 9456 19252 9462 19264
rect 7834 19184 7840 19236
rect 7892 19224 7898 19236
rect 10778 19224 10784 19236
rect 7892 19196 10784 19224
rect 7892 19184 7898 19196
rect 10778 19184 10784 19196
rect 10836 19184 10842 19236
rect 11241 19227 11299 19233
rect 11241 19193 11253 19227
rect 11287 19224 11299 19227
rect 11422 19224 11428 19236
rect 11287 19196 11428 19224
rect 11287 19193 11299 19196
rect 11241 19187 11299 19193
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 14642 19184 14648 19236
rect 14700 19224 14706 19236
rect 15933 19227 15991 19233
rect 15933 19224 15945 19227
rect 14700 19196 15945 19224
rect 14700 19184 14706 19196
rect 15933 19193 15945 19196
rect 15979 19193 15991 19227
rect 16500 19224 16528 19264
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16632 19264 16957 19292
rect 16632 19252 16638 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 21634 19292 21640 19304
rect 20763 19264 21640 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 22833 19295 22891 19301
rect 22833 19261 22845 19295
rect 22879 19292 22891 19295
rect 23290 19292 23296 19304
rect 22879 19264 23296 19292
rect 22879 19261 22891 19264
rect 22833 19255 22891 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 18782 19224 18788 19236
rect 16500 19196 18788 19224
rect 15933 19187 15991 19193
rect 18782 19184 18788 19196
rect 18840 19184 18846 19236
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 9582 19156 9588 19168
rect 8352 19128 9588 19156
rect 8352 19116 8358 19128
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14458 19156 14464 19168
rect 13964 19128 14464 19156
rect 13964 19116 13970 19128
rect 14458 19116 14464 19128
rect 14516 19156 14522 19168
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 14516 19128 14565 19156
rect 14516 19116 14522 19128
rect 14553 19125 14565 19128
rect 14599 19156 14611 19159
rect 15102 19156 15108 19168
rect 14599 19128 15108 19156
rect 14599 19125 14611 19128
rect 14553 19119 14611 19125
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 19150 19116 19156 19168
rect 19208 19116 19214 19168
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 21818 19116 21824 19168
rect 21876 19116 21882 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 8389 18955 8447 18961
rect 8389 18921 8401 18955
rect 8435 18952 8447 18955
rect 8478 18952 8484 18964
rect 8435 18924 8484 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 8478 18912 8484 18924
rect 8536 18952 8542 18964
rect 9306 18952 9312 18964
rect 8536 18924 9312 18952
rect 8536 18912 8542 18924
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 10781 18955 10839 18961
rect 10781 18921 10793 18955
rect 10827 18952 10839 18955
rect 10870 18952 10876 18964
rect 10827 18924 10876 18952
rect 10827 18921 10839 18924
rect 10781 18915 10839 18921
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 12253 18955 12311 18961
rect 12253 18921 12265 18955
rect 12299 18952 12311 18955
rect 14550 18952 14556 18964
rect 12299 18924 14556 18952
rect 12299 18921 12311 18924
rect 12253 18915 12311 18921
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 17552 18924 17877 18952
rect 17552 18912 17558 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 17865 18915 17923 18921
rect 25225 18955 25283 18961
rect 25225 18921 25237 18955
rect 25271 18952 25283 18955
rect 26786 18952 26792 18964
rect 25271 18924 26792 18952
rect 25271 18921 25283 18924
rect 25225 18915 25283 18921
rect 10042 18844 10048 18896
rect 10100 18884 10106 18896
rect 12713 18887 12771 18893
rect 12713 18884 12725 18887
rect 10100 18856 12725 18884
rect 10100 18844 10106 18856
rect 12713 18853 12725 18856
rect 12759 18853 12771 18887
rect 12713 18847 12771 18853
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8294 18816 8300 18828
rect 6963 18788 8300 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 10502 18816 10508 18828
rect 10275 18788 10508 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 11020 18788 11621 18816
rect 11020 18776 11026 18788
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 11793 18819 11851 18825
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 12618 18816 12624 18828
rect 11839 18788 12624 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 13265 18819 13323 18825
rect 13265 18785 13277 18819
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6604 18720 6653 18748
rect 6604 18708 6610 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 13280 18748 13308 18779
rect 16390 18776 16396 18828
rect 16448 18816 16454 18828
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16448 18788 16957 18816
rect 16448 18776 16454 18788
rect 16945 18785 16957 18788
rect 16991 18785 17003 18819
rect 16945 18779 17003 18785
rect 19150 18776 19156 18828
rect 19208 18816 19214 18828
rect 19208 18788 22048 18816
rect 19208 18776 19214 18788
rect 10836 18720 13308 18748
rect 17221 18751 17279 18757
rect 10836 18708 10842 18720
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17494 18748 17500 18760
rect 17267 18720 17500 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 22020 18757 22048 18788
rect 23842 18776 23848 18828
rect 23900 18776 23906 18828
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 8294 18680 8300 18692
rect 8142 18652 8300 18680
rect 8294 18640 8300 18652
rect 8352 18680 8358 18692
rect 8665 18683 8723 18689
rect 8665 18680 8677 18683
rect 8352 18652 8677 18680
rect 8352 18640 8358 18652
rect 8665 18649 8677 18652
rect 8711 18649 8723 18683
rect 8665 18643 8723 18649
rect 8846 18640 8852 18692
rect 8904 18680 8910 18692
rect 9398 18680 9404 18692
rect 8904 18652 9404 18680
rect 8904 18640 8910 18652
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 10413 18683 10471 18689
rect 10413 18680 10425 18683
rect 9692 18652 10425 18680
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 9214 18612 9220 18624
rect 8812 18584 9220 18612
rect 8812 18572 8818 18584
rect 9214 18572 9220 18584
rect 9272 18612 9278 18624
rect 9692 18621 9720 18652
rect 10413 18649 10425 18652
rect 10459 18649 10471 18683
rect 10413 18643 10471 18649
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 11057 18683 11115 18689
rect 11057 18680 11069 18683
rect 10560 18652 11069 18680
rect 10560 18640 10566 18652
rect 11057 18649 11069 18652
rect 11103 18649 11115 18683
rect 11057 18643 11115 18649
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9272 18584 9689 18612
rect 9272 18572 9278 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9677 18575 9735 18581
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 11072 18612 11100 18643
rect 11146 18640 11152 18692
rect 11204 18680 11210 18692
rect 11885 18683 11943 18689
rect 11885 18680 11897 18683
rect 11204 18652 11897 18680
rect 11204 18640 11210 18652
rect 11885 18649 11897 18652
rect 11931 18649 11943 18683
rect 17678 18680 17684 18692
rect 11885 18643 11943 18649
rect 17236 18652 17684 18680
rect 17236 18624 17264 18652
rect 17678 18640 17684 18652
rect 17736 18680 17742 18692
rect 18049 18683 18107 18689
rect 18049 18680 18061 18683
rect 17736 18652 18061 18680
rect 17736 18640 17742 18652
rect 18049 18649 18061 18652
rect 18095 18649 18107 18683
rect 21468 18680 21496 18711
rect 22738 18708 22744 18760
rect 22796 18708 22802 18760
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18748 24823 18751
rect 25240 18748 25268 18915
rect 26786 18912 26792 18924
rect 26844 18912 26850 18964
rect 24811 18720 25268 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 24486 18680 24492 18692
rect 21468 18652 24492 18680
rect 18049 18643 18107 18649
rect 24486 18640 24492 18652
rect 24544 18640 24550 18692
rect 11514 18612 11520 18624
rect 11072 18584 11520 18612
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12860 18584 13093 18612
rect 12860 18572 12866 18584
rect 13081 18581 13093 18584
rect 13127 18581 13139 18615
rect 13081 18575 13139 18581
rect 13173 18615 13231 18621
rect 13173 18581 13185 18615
rect 13219 18612 13231 18615
rect 13262 18612 13268 18624
rect 13219 18584 13268 18612
rect 13219 18581 13231 18584
rect 13173 18575 13231 18581
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13817 18615 13875 18621
rect 13817 18581 13829 18615
rect 13863 18612 13875 18615
rect 14182 18612 14188 18624
rect 13863 18584 14188 18612
rect 13863 18581 13875 18584
rect 13817 18575 13875 18581
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 14274 18572 14280 18624
rect 14332 18572 14338 18624
rect 17129 18615 17187 18621
rect 17129 18581 17141 18615
rect 17175 18612 17187 18615
rect 17218 18612 17224 18624
rect 17175 18584 17224 18612
rect 17175 18581 17187 18584
rect 17129 18575 17187 18581
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 17589 18615 17647 18621
rect 17589 18612 17601 18615
rect 17552 18584 17601 18612
rect 17552 18572 17558 18584
rect 17589 18581 17601 18584
rect 17635 18581 17647 18615
rect 17589 18575 17647 18581
rect 20898 18572 20904 18624
rect 20956 18612 20962 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 20956 18584 21281 18612
rect 20956 18572 20962 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 22186 18572 22192 18624
rect 22244 18572 22250 18624
rect 24670 18572 24676 18624
rect 24728 18572 24734 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 6546 18368 6552 18420
rect 6604 18408 6610 18420
rect 9122 18408 9128 18420
rect 6604 18380 9128 18408
rect 6604 18368 6610 18380
rect 9122 18368 9128 18380
rect 9180 18408 9186 18420
rect 9180 18380 9536 18408
rect 9180 18368 9186 18380
rect 8202 18300 8208 18352
rect 8260 18300 8266 18352
rect 9508 18284 9536 18380
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 10376 18380 13829 18408
rect 10376 18368 10382 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 14240 18380 14289 18408
rect 14240 18368 14246 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14921 18411 14979 18417
rect 14921 18377 14933 18411
rect 14967 18408 14979 18411
rect 16574 18408 16580 18420
rect 14967 18380 16580 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 10229 18343 10287 18349
rect 10229 18309 10241 18343
rect 10275 18340 10287 18343
rect 11238 18340 11244 18352
rect 10275 18312 11244 18340
rect 10275 18309 10287 18312
rect 10229 18303 10287 18309
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 12066 18340 12072 18352
rect 11532 18312 12072 18340
rect 9490 18232 9496 18284
rect 9548 18232 9554 18284
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10321 18275 10379 18281
rect 9640 18244 10088 18272
rect 9640 18232 9646 18244
rect 7742 18164 7748 18216
rect 7800 18164 7806 18216
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 9674 18204 9680 18216
rect 9263 18176 9680 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 10060 18213 10088 18244
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 11057 18275 11115 18281
rect 11057 18241 11069 18275
rect 11103 18272 11115 18275
rect 11330 18272 11336 18284
rect 11103 18244 11336 18272
rect 11103 18241 11115 18244
rect 11057 18235 11115 18241
rect 10045 18207 10103 18213
rect 10045 18173 10057 18207
rect 10091 18173 10103 18207
rect 10045 18167 10103 18173
rect 7558 18028 7564 18080
rect 7616 18068 7622 18080
rect 10336 18068 10364 18235
rect 11330 18232 11336 18244
rect 11388 18272 11394 18284
rect 11532 18272 11560 18312
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 13265 18343 13323 18349
rect 13265 18309 13277 18343
rect 13311 18340 13323 18343
rect 13354 18340 13360 18352
rect 13311 18312 13360 18340
rect 13311 18309 13323 18312
rect 13265 18303 13323 18309
rect 13354 18300 13360 18312
rect 13412 18300 13418 18352
rect 11388 18244 11560 18272
rect 11388 18232 11394 18244
rect 11606 18232 11612 18284
rect 11664 18272 11670 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 11664 18244 12449 18272
rect 11664 18232 11670 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18272 14243 18275
rect 14936 18272 14964 18371
rect 16574 18368 16580 18380
rect 16632 18408 16638 18420
rect 25866 18408 25872 18420
rect 16632 18380 25872 18408
rect 16632 18368 16638 18380
rect 25866 18368 25872 18380
rect 25924 18368 25930 18420
rect 23293 18343 23351 18349
rect 23293 18309 23305 18343
rect 23339 18340 23351 18343
rect 24854 18340 24860 18352
rect 23339 18312 24860 18340
rect 23339 18309 23351 18312
rect 23293 18303 23351 18309
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 14231 18244 14964 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 18262 18244 19012 18272
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 11882 18204 11888 18216
rect 11296 18176 11888 18204
rect 11296 18164 11302 18176
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 13504 18176 14381 18204
rect 13504 18164 13510 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 16816 18176 17141 18204
rect 16816 18164 16822 18176
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 15010 18136 15016 18148
rect 10735 18108 15016 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 15010 18096 15016 18108
rect 15068 18096 15074 18148
rect 16960 18080 16988 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17129 18167 17187 18173
rect 7616 18040 10364 18068
rect 7616 18028 7622 18040
rect 16942 18028 16948 18080
rect 17000 18028 17006 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18984 18077 19012 18244
rect 21266 18232 21272 18284
rect 21324 18232 21330 18284
rect 22186 18232 22192 18284
rect 22244 18232 22250 18284
rect 23474 18232 23480 18284
rect 23532 18272 23538 18284
rect 23937 18275 23995 18281
rect 23937 18272 23949 18275
rect 23532 18244 23949 18272
rect 23532 18232 23538 18244
rect 23937 18241 23949 18244
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 24578 18164 24584 18216
rect 24636 18164 24642 18216
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 18380 18040 18613 18068
rect 18380 18028 18386 18040
rect 18601 18037 18613 18040
rect 18647 18037 18659 18071
rect 18601 18031 18659 18037
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19150 18068 19156 18080
rect 19015 18040 19156 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 21082 18028 21088 18080
rect 21140 18028 21146 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 8570 17824 8576 17876
rect 8628 17824 8634 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 11238 17864 11244 17876
rect 9732 17836 11244 17864
rect 9732 17824 9738 17836
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13998 17864 14004 17876
rect 13035 17836 14004 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 17920 17836 18429 17864
rect 17920 17824 17926 17836
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 24854 17864 24860 17876
rect 18417 17827 18475 17833
rect 23308 17836 24860 17864
rect 13446 17796 13452 17808
rect 12268 17768 13452 17796
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7892 17700 7941 17728
rect 7892 17688 7898 17700
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 9490 17688 9496 17740
rect 9548 17728 9554 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 9548 17700 9781 17728
rect 9548 17688 9554 17700
rect 9769 17697 9781 17700
rect 9815 17697 9827 17731
rect 9769 17691 9827 17697
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10134 17728 10140 17740
rect 10091 17700 10140 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10134 17688 10140 17700
rect 10192 17728 10198 17740
rect 12268 17728 12296 17768
rect 13446 17756 13452 17768
rect 13504 17756 13510 17808
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 14185 17799 14243 17805
rect 14185 17796 14197 17799
rect 13872 17768 14197 17796
rect 13872 17756 13878 17768
rect 14185 17765 14197 17768
rect 14231 17796 14243 17799
rect 16666 17796 16672 17808
rect 14231 17768 16672 17796
rect 14231 17765 14243 17768
rect 14185 17759 14243 17765
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 21453 17799 21511 17805
rect 21453 17765 21465 17799
rect 21499 17796 21511 17799
rect 23198 17796 23204 17808
rect 21499 17768 23204 17796
rect 21499 17765 21511 17768
rect 21453 17759 21511 17765
rect 23198 17756 23204 17768
rect 23256 17756 23262 17808
rect 10192 17700 12296 17728
rect 12437 17731 12495 17737
rect 10192 17688 10198 17700
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 12526 17728 12532 17740
rect 12483 17700 12532 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 17310 17728 17316 17740
rect 16991 17700 17316 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 17678 17688 17684 17740
rect 17736 17728 17742 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17736 17700 17969 17728
rect 17736 17688 17742 17700
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 23308 17737 23336 17836
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 26142 17796 26148 17808
rect 24044 17768 26148 17796
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 18380 17700 19533 17728
rect 18380 17688 18386 17700
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 23293 17731 23351 17737
rect 23293 17697 23305 17731
rect 23339 17697 23351 17731
rect 24044 17728 24072 17768
rect 26142 17756 26148 17768
rect 26200 17756 26206 17808
rect 23293 17691 23351 17697
rect 23492 17700 24072 17728
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17660 8171 17663
rect 8159 17632 9812 17660
rect 8159 17629 8171 17632
rect 8113 17623 8171 17629
rect 7650 17552 7656 17604
rect 7708 17592 7714 17604
rect 8205 17595 8263 17601
rect 8205 17592 8217 17595
rect 7708 17564 8217 17592
rect 7708 17552 7714 17564
rect 8205 17561 8217 17564
rect 8251 17561 8263 17595
rect 8205 17555 8263 17561
rect 7374 17484 7380 17536
rect 7432 17484 7438 17536
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9398 17524 9404 17536
rect 9355 17496 9404 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9784 17524 9812 17632
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11572 17632 11805 17660
rect 11572 17620 11578 17632
rect 11793 17629 11805 17632
rect 11839 17660 11851 17663
rect 11882 17660 11888 17672
rect 11839 17632 11888 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 14274 17660 14280 17672
rect 12667 17632 14280 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16758 17660 16764 17672
rect 16715 17632 16764 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 17773 17663 17831 17669
rect 17773 17660 17785 17663
rect 17644 17632 17785 17660
rect 17644 17620 17650 17632
rect 17773 17629 17785 17632
rect 17819 17660 17831 17663
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 17819 17632 18797 17660
rect 17819 17629 17831 17632
rect 17773 17623 17831 17629
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19484 17632 19717 17660
rect 19484 17620 19490 17632
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 11330 17592 11336 17604
rect 11270 17564 11336 17592
rect 11330 17552 11336 17564
rect 11388 17592 11394 17604
rect 11974 17592 11980 17604
rect 11388 17564 11980 17592
rect 11388 17552 11394 17564
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 12529 17595 12587 17601
rect 12529 17592 12541 17595
rect 12406 17564 12541 17592
rect 10226 17524 10232 17536
rect 9784 17496 10232 17524
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 12406 17524 12434 17564
rect 12529 17561 12541 17564
rect 12575 17592 12587 17595
rect 14182 17592 14188 17604
rect 12575 17564 14188 17592
rect 12575 17561 12587 17564
rect 12529 17555 12587 17561
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 16356 17564 18736 17592
rect 16356 17552 16362 17564
rect 12124 17496 12434 17524
rect 12124 17484 12130 17496
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13228 17496 13461 17524
rect 13228 17484 13234 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 13449 17487 13507 17493
rect 15654 17484 15660 17536
rect 15712 17484 15718 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 17184 17496 17417 17524
rect 17184 17484 17190 17496
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 17405 17487 17463 17493
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 17828 17496 17877 17524
rect 17828 17484 17834 17496
rect 17865 17493 17877 17496
rect 17911 17524 17923 17527
rect 18414 17524 18420 17536
rect 17911 17496 18420 17524
rect 17911 17493 17923 17496
rect 17865 17487 17923 17493
rect 18414 17484 18420 17496
rect 18472 17524 18478 17536
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 18472 17496 18613 17524
rect 18472 17484 18478 17496
rect 18601 17493 18613 17496
rect 18647 17493 18659 17527
rect 18708 17524 18736 17564
rect 19242 17552 19248 17604
rect 19300 17592 19306 17604
rect 20640 17592 20668 17623
rect 21174 17620 21180 17672
rect 21232 17660 21238 17672
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 21232 17632 21281 17660
rect 21232 17620 21238 17632
rect 21269 17629 21281 17632
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 21910 17620 21916 17672
rect 21968 17620 21974 17672
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17660 22155 17663
rect 22186 17660 22192 17672
rect 22143 17632 22192 17660
rect 22143 17629 22155 17632
rect 22097 17623 22155 17629
rect 22186 17620 22192 17632
rect 22244 17660 22250 17672
rect 23492 17660 23520 17700
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 22244 17632 23520 17660
rect 22244 17620 22250 17632
rect 23658 17620 23664 17672
rect 23716 17660 23722 17672
rect 23845 17663 23903 17669
rect 23845 17660 23857 17663
rect 23716 17632 23857 17660
rect 23716 17620 23722 17632
rect 23845 17629 23857 17632
rect 23891 17629 23903 17663
rect 23845 17623 23903 17629
rect 24394 17592 24400 17604
rect 19300 17564 20668 17592
rect 20824 17564 22094 17592
rect 19300 17552 19306 17564
rect 19797 17527 19855 17533
rect 19797 17524 19809 17527
rect 18708 17496 19809 17524
rect 18601 17487 18659 17493
rect 19797 17493 19809 17496
rect 19843 17493 19855 17527
rect 19797 17487 19855 17493
rect 20165 17527 20223 17533
rect 20165 17493 20177 17527
rect 20211 17524 20223 17527
rect 20714 17524 20720 17536
rect 20211 17496 20720 17524
rect 20211 17493 20223 17496
rect 20165 17487 20223 17493
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 20824 17533 20852 17564
rect 20809 17527 20867 17533
rect 20809 17493 20821 17527
rect 20855 17493 20867 17527
rect 22066 17524 22094 17564
rect 22296 17564 24400 17592
rect 22296 17524 22324 17564
rect 24394 17552 24400 17564
rect 24452 17552 24458 17604
rect 22066 17496 22324 17524
rect 20809 17487 20867 17493
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 22612 17496 24593 17524
rect 22612 17484 22618 17496
rect 24581 17493 24593 17496
rect 24627 17493 24639 17527
rect 24581 17487 24639 17493
rect 24762 17484 24768 17536
rect 24820 17524 24826 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24820 17496 24961 17524
rect 24820 17484 24826 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7432 17292 8033 17320
rect 7432 17280 7438 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 9769 17323 9827 17329
rect 9769 17289 9781 17323
rect 9815 17320 9827 17323
rect 11054 17320 11060 17332
rect 9815 17292 11060 17320
rect 9815 17289 9827 17292
rect 9769 17283 9827 17289
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11330 17320 11336 17332
rect 11164 17292 11336 17320
rect 9490 17212 9496 17264
rect 9548 17252 9554 17264
rect 11164 17261 11192 17292
rect 11330 17280 11336 17292
rect 11388 17320 11394 17332
rect 11606 17320 11612 17332
rect 11388 17292 11612 17320
rect 11388 17280 11394 17292
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12250 17320 12256 17332
rect 12032 17292 12256 17320
rect 12032 17280 12038 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 13170 17280 13176 17332
rect 13228 17280 13234 17332
rect 13541 17323 13599 17329
rect 13541 17289 13553 17323
rect 13587 17320 13599 17323
rect 15378 17320 15384 17332
rect 13587 17292 15384 17320
rect 13587 17289 13599 17292
rect 13541 17283 13599 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15746 17320 15752 17332
rect 15672 17292 15752 17320
rect 10321 17255 10379 17261
rect 10321 17252 10333 17255
rect 9548 17224 10333 17252
rect 9548 17212 9554 17224
rect 10321 17221 10333 17224
rect 10367 17221 10379 17255
rect 10321 17215 10379 17221
rect 11149 17255 11207 17261
rect 11149 17221 11161 17255
rect 11195 17221 11207 17255
rect 15672 17252 15700 17292
rect 15746 17280 15752 17292
rect 15804 17320 15810 17332
rect 17310 17320 17316 17332
rect 15804 17292 17316 17320
rect 15804 17280 15810 17292
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 20220 17292 20361 17320
rect 20220 17280 20226 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 22005 17323 22063 17329
rect 22005 17289 22017 17323
rect 22051 17320 22063 17323
rect 22186 17320 22192 17332
rect 22051 17292 22192 17320
rect 22051 17289 22063 17292
rect 22005 17283 22063 17289
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22741 17323 22799 17329
rect 22741 17289 22753 17323
rect 22787 17320 22799 17323
rect 24118 17320 24124 17332
rect 22787 17292 24124 17320
rect 22787 17289 22799 17292
rect 22741 17283 22799 17289
rect 24118 17280 24124 17292
rect 24176 17280 24182 17332
rect 15594 17224 15700 17252
rect 11149 17215 11207 17221
rect 15930 17212 15936 17264
rect 15988 17252 15994 17264
rect 17037 17255 17095 17261
rect 15988 17224 16988 17252
rect 15988 17212 15994 17224
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7432 17156 7941 17184
rect 7432 17144 7438 17156
rect 7929 17153 7941 17156
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 8938 17184 8944 17196
rect 8803 17156 8944 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 8938 17144 8944 17156
rect 8996 17184 9002 17196
rect 9309 17187 9367 17193
rect 9309 17184 9321 17187
rect 8996 17156 9321 17184
rect 8996 17144 9002 17156
rect 9309 17153 9321 17156
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16850 17184 16856 17196
rect 16347 17156 16856 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 16960 17184 16988 17224
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 17862 17252 17868 17264
rect 17083 17224 17868 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 18049 17255 18107 17261
rect 18049 17221 18061 17255
rect 18095 17252 18107 17255
rect 18506 17252 18512 17264
rect 18095 17224 18512 17252
rect 18095 17221 18107 17224
rect 18049 17215 18107 17221
rect 18506 17212 18512 17224
rect 18564 17212 18570 17264
rect 18782 17212 18788 17264
rect 18840 17252 18846 17264
rect 18877 17255 18935 17261
rect 18877 17252 18889 17255
rect 18840 17224 18889 17252
rect 18840 17212 18846 17224
rect 18877 17221 18889 17224
rect 18923 17221 18935 17255
rect 20625 17255 20683 17261
rect 20625 17252 20637 17255
rect 20102 17224 20637 17252
rect 18877 17215 18935 17221
rect 20625 17221 20637 17224
rect 20671 17252 20683 17255
rect 20990 17252 20996 17264
rect 20671 17224 20996 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 20990 17212 20996 17224
rect 21048 17252 21054 17264
rect 21818 17252 21824 17264
rect 21048 17224 21824 17252
rect 21048 17212 21054 17224
rect 21818 17212 21824 17224
rect 21876 17252 21882 17264
rect 22278 17252 22284 17264
rect 21876 17224 22284 17252
rect 21876 17212 21882 17224
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 23750 17212 23756 17264
rect 23808 17212 23814 17264
rect 24026 17212 24032 17264
rect 24084 17252 24090 17264
rect 24084 17224 24242 17252
rect 24084 17212 24090 17224
rect 21453 17187 21511 17193
rect 16960 17156 17908 17184
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17116 7895 17119
rect 8386 17116 8392 17128
rect 7883 17088 8392 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 9214 17076 9220 17128
rect 9272 17076 9278 17128
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12768 17088 12909 17116
rect 12768 17076 12774 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13630 17116 13636 17128
rect 13127 17088 13636 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 11514 17008 11520 17060
rect 11572 17048 11578 17060
rect 12066 17048 12072 17060
rect 11572 17020 12072 17048
rect 11572 17008 11578 17020
rect 12066 17008 12072 17020
rect 12124 17008 12130 17060
rect 12529 17051 12587 17057
rect 12529 17017 12541 17051
rect 12575 17048 12587 17051
rect 13096 17048 13124 17079
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 14826 17116 14832 17128
rect 14608 17088 14832 17116
rect 14608 17076 14614 17088
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 16022 17076 16028 17128
rect 16080 17076 16086 17128
rect 17880 17125 17908 17156
rect 21453 17153 21465 17187
rect 21499 17184 21511 17187
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 21499 17156 22661 17184
rect 21499 17153 21511 17156
rect 21453 17147 21511 17153
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 18598 17076 18604 17128
rect 18656 17076 18662 17128
rect 22925 17119 22983 17125
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 22971 17088 25237 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 25225 17085 25237 17088
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 12575 17020 13124 17048
rect 12575 17017 12587 17020
rect 12529 17011 12587 17017
rect 20438 17008 20444 17060
rect 20496 17048 20502 17060
rect 22940 17048 22968 17079
rect 20496 17020 22968 17048
rect 20496 17008 20502 17020
rect 8389 16983 8447 16989
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 11790 16980 11796 16992
rect 8435 16952 11796 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16264 16952 16957 16980
rect 16264 16940 16270 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 17497 16983 17555 16989
rect 17497 16949 17509 16983
rect 17543 16980 17555 16983
rect 17586 16980 17592 16992
rect 17543 16952 17592 16980
rect 17543 16949 17555 16952
rect 17497 16943 17555 16949
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 22281 16983 22339 16989
rect 22281 16949 22293 16983
rect 22327 16980 22339 16983
rect 22370 16980 22376 16992
rect 22327 16952 22376 16980
rect 22327 16949 22339 16952
rect 22281 16943 22339 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23198 16940 23204 16992
rect 23256 16980 23262 16992
rect 23934 16980 23940 16992
rect 23256 16952 23940 16980
rect 23256 16940 23262 16952
rect 23934 16940 23940 16952
rect 23992 16940 23998 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 8444 16748 8493 16776
rect 8444 16736 8450 16748
rect 8481 16745 8493 16748
rect 8527 16745 8539 16779
rect 13262 16776 13268 16788
rect 8481 16739 8539 16745
rect 11900 16748 13268 16776
rect 11238 16708 11244 16720
rect 10428 16680 11244 16708
rect 10428 16649 10456 16680
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 11900 16640 11928 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 13909 16779 13967 16785
rect 13909 16745 13921 16779
rect 13955 16776 13967 16779
rect 14458 16776 14464 16788
rect 13955 16748 14464 16776
rect 13955 16745 13967 16748
rect 13909 16739 13967 16745
rect 13924 16708 13952 16739
rect 14458 16736 14464 16748
rect 14516 16776 14522 16788
rect 15746 16776 15752 16788
rect 14516 16748 15752 16776
rect 14516 16736 14522 16748
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 21266 16776 21272 16788
rect 20180 16748 21272 16776
rect 13648 16680 13952 16708
rect 10551 16612 11928 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 13170 16640 13176 16652
rect 12584 16612 13176 16640
rect 12584 16600 12590 16612
rect 13170 16600 13176 16612
rect 13228 16640 13234 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 13228 16612 13277 16640
rect 13228 16600 13234 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 13538 16600 13544 16652
rect 13596 16600 13602 16652
rect 13648 16572 13676 16680
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 13556 16544 13676 16572
rect 13740 16612 14657 16640
rect 10410 16464 10416 16516
rect 10468 16504 10474 16516
rect 13556 16504 13584 16544
rect 10468 16476 11008 16504
rect 12834 16476 13584 16504
rect 10468 16464 10474 16476
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 10594 16436 10600 16448
rect 9916 16408 10600 16436
rect 9916 16396 9922 16408
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 10980 16445 11008 16476
rect 10965 16439 11023 16445
rect 10965 16405 10977 16439
rect 11011 16405 11023 16439
rect 10965 16399 11023 16405
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 13740 16436 13768 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 15838 16600 15844 16652
rect 15896 16600 15902 16652
rect 16850 16600 16856 16652
rect 16908 16640 16914 16652
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 16908 16612 17969 16640
rect 16908 16600 16914 16612
rect 17957 16609 17969 16612
rect 18003 16640 18015 16643
rect 18598 16640 18604 16652
rect 18003 16612 18604 16640
rect 18003 16609 18015 16612
rect 17957 16603 18015 16609
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 15654 16532 15660 16584
rect 15712 16572 15718 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15712 16544 16129 16572
rect 15712 16532 15718 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 16117 16535 16175 16541
rect 16592 16544 18705 16572
rect 16592 16504 16620 16544
rect 18693 16541 18705 16544
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20180 16572 20208 16748
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22738 16776 22744 16788
rect 22336 16748 22744 16776
rect 22336 16736 22342 16748
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 24581 16779 24639 16785
rect 24581 16776 24593 16779
rect 23716 16748 24593 16776
rect 23716 16736 23722 16748
rect 24581 16745 24593 16748
rect 24627 16745 24639 16779
rect 24581 16739 24639 16745
rect 20254 16600 20260 16652
rect 20312 16600 20318 16652
rect 20530 16600 20536 16652
rect 20588 16600 20594 16652
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 20680 16612 22017 16640
rect 20680 16600 20686 16612
rect 19843 16544 20208 16572
rect 21928 16572 21956 16612
rect 22005 16609 22017 16612
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 22278 16572 22284 16584
rect 21928 16544 22284 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 23842 16532 23848 16584
rect 23900 16532 23906 16584
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 15304 16476 16620 16504
rect 11848 16408 13768 16436
rect 11848 16396 11854 16408
rect 14182 16396 14188 16448
rect 14240 16396 14246 16448
rect 14826 16396 14832 16448
rect 14884 16396 14890 16448
rect 14918 16396 14924 16448
rect 14976 16396 14982 16448
rect 15304 16445 15332 16476
rect 16666 16464 16672 16516
rect 16724 16504 16730 16516
rect 17221 16507 17279 16513
rect 17221 16504 17233 16507
rect 16724 16476 17233 16504
rect 16724 16464 16730 16476
rect 17221 16473 17233 16476
rect 17267 16504 17279 16507
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 17267 16476 19257 16504
rect 17267 16473 17279 16476
rect 17221 16467 17279 16473
rect 19245 16473 19257 16476
rect 19291 16504 19303 16507
rect 19334 16504 19340 16516
rect 19291 16476 19340 16504
rect 19291 16473 19303 16476
rect 19245 16467 19303 16473
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 19444 16476 20484 16504
rect 15289 16439 15347 16445
rect 15289 16405 15301 16439
rect 15335 16405 15347 16439
rect 15289 16399 15347 16405
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 16114 16436 16120 16448
rect 16071 16408 16120 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 16482 16396 16488 16448
rect 16540 16396 16546 16448
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 17310 16436 17316 16448
rect 16908 16408 17316 16436
rect 16908 16396 16914 16408
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 18877 16439 18935 16445
rect 18877 16405 18889 16439
rect 18923 16436 18935 16439
rect 19444 16436 19472 16476
rect 18923 16408 19472 16436
rect 18923 16405 18935 16408
rect 18877 16399 18935 16405
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19613 16439 19671 16445
rect 19613 16436 19625 16439
rect 19576 16408 19625 16436
rect 19576 16396 19582 16408
rect 19613 16405 19625 16408
rect 19659 16405 19671 16439
rect 20456 16436 20484 16476
rect 20990 16464 20996 16516
rect 21048 16464 21054 16516
rect 24780 16504 24808 16535
rect 21836 16476 24808 16504
rect 21836 16436 21864 16476
rect 20456 16408 21864 16436
rect 19613 16399 19671 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 11882 16192 11888 16244
rect 11940 16192 11946 16244
rect 12158 16192 12164 16244
rect 12216 16192 12222 16244
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13357 16235 13415 16241
rect 13357 16232 13369 16235
rect 13320 16204 13369 16232
rect 13320 16192 13326 16204
rect 13357 16201 13369 16204
rect 13403 16201 13415 16235
rect 13357 16195 13415 16201
rect 13725 16235 13783 16241
rect 13725 16201 13737 16235
rect 13771 16232 13783 16235
rect 14182 16232 14188 16244
rect 13771 16204 14188 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 14826 16232 14832 16244
rect 14599 16204 14832 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 14976 16204 15761 16232
rect 14976 16192 14982 16204
rect 15749 16201 15761 16204
rect 15795 16201 15807 16235
rect 15749 16195 15807 16201
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16724 16204 16773 16232
rect 16724 16192 16730 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 19978 16232 19984 16244
rect 16761 16195 16819 16201
rect 19904 16204 19984 16232
rect 8294 16164 8300 16176
rect 8050 16136 8300 16164
rect 8294 16124 8300 16136
rect 8352 16164 8358 16176
rect 8570 16164 8576 16176
rect 8352 16136 8576 16164
rect 8352 16124 8358 16136
rect 8570 16124 8576 16136
rect 8628 16124 8634 16176
rect 11330 16124 11336 16176
rect 11388 16164 11394 16176
rect 13814 16164 13820 16176
rect 11388 16136 13820 16164
rect 11388 16124 11394 16136
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 14200 16164 14228 16192
rect 14200 16136 17264 16164
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13998 16096 14004 16108
rect 12575 16068 14004 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 17236 16096 17264 16136
rect 17310 16124 17316 16176
rect 17368 16124 17374 16176
rect 18874 16164 18880 16176
rect 18064 16136 18880 16164
rect 17954 16096 17960 16108
rect 17236 16068 17960 16096
rect 14921 16059 14979 16065
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18064 16105 18092 16136
rect 18874 16124 18880 16136
rect 18932 16124 18938 16176
rect 19245 16167 19303 16173
rect 19245 16133 19257 16167
rect 19291 16164 19303 16167
rect 19334 16164 19340 16176
rect 19291 16136 19340 16164
rect 19291 16133 19303 16136
rect 19245 16127 19303 16133
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19904 16096 19932 16204
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 20254 16232 20260 16244
rect 20088 16204 20260 16232
rect 20088 16173 20116 16204
rect 20254 16192 20260 16204
rect 20312 16232 20318 16244
rect 23566 16232 23572 16244
rect 20312 16204 23572 16232
rect 20312 16192 20318 16204
rect 20073 16167 20131 16173
rect 20073 16133 20085 16167
rect 20119 16133 20131 16167
rect 20073 16127 20131 16133
rect 20346 16124 20352 16176
rect 20404 16164 20410 16176
rect 20993 16167 21051 16173
rect 20993 16164 21005 16167
rect 20404 16136 21005 16164
rect 20404 16124 20410 16136
rect 20993 16133 21005 16136
rect 21039 16133 21051 16167
rect 20993 16127 21051 16133
rect 18739 16068 19932 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 22020 16105 22048 16204
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 22278 16124 22284 16176
rect 22336 16124 22342 16176
rect 22738 16124 22744 16176
rect 22796 16124 22802 16176
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20036 16068 21097 16096
rect 20036 16056 20042 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 23900 16068 24777 16096
rect 23900 16056 23906 16068
rect 24765 16065 24777 16068
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 6822 15988 6828 16040
rect 6880 15988 6886 16040
rect 12618 15988 12624 16040
rect 12676 15988 12682 16040
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 8662 15960 8668 15972
rect 8312 15932 8668 15960
rect 8312 15904 8340 15932
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 11882 15920 11888 15972
rect 11940 15960 11946 15972
rect 12728 15960 12756 15991
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13688 16000 13829 16028
rect 13688 15988 13694 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 11940 15932 12756 15960
rect 11940 15920 11946 15932
rect 13446 15920 13452 15972
rect 13504 15960 13510 15972
rect 13924 15960 13952 15991
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 15997 15163 16031
rect 15105 15991 15163 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 13504 15932 13952 15960
rect 13504 15920 13510 15932
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 8570 15852 8576 15904
rect 8628 15852 8634 15904
rect 13170 15852 13176 15904
rect 13228 15892 13234 15904
rect 15120 15892 15148 15991
rect 16574 15920 16580 15972
rect 16632 15960 16638 15972
rect 17865 15963 17923 15969
rect 17865 15960 17877 15963
rect 16632 15932 17877 15960
rect 16632 15920 16638 15932
rect 17865 15929 17877 15932
rect 17911 15929 17923 15963
rect 20916 15960 20944 15991
rect 22738 15988 22744 16040
rect 22796 16028 22802 16040
rect 24026 16028 24032 16040
rect 22796 16000 24032 16028
rect 22796 15988 22802 16000
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24489 16031 24547 16037
rect 24489 15997 24501 16031
rect 24535 16028 24547 16031
rect 24578 16028 24584 16040
rect 24535 16000 24584 16028
rect 24535 15997 24547 16000
rect 24489 15991 24547 15997
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 20916 15932 22094 15960
rect 17865 15923 17923 15929
rect 13228 15864 15148 15892
rect 13228 15852 13234 15864
rect 16114 15852 16120 15904
rect 16172 15892 16178 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 16172 15864 16221 15892
rect 16172 15852 16178 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16209 15855 16267 15861
rect 17218 15852 17224 15904
rect 17276 15852 17282 15904
rect 18509 15895 18567 15901
rect 18509 15861 18521 15895
rect 18555 15892 18567 15895
rect 19242 15892 19248 15904
rect 18555 15864 19248 15892
rect 18555 15861 18567 15864
rect 18509 15855 18567 15861
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 21450 15852 21456 15904
rect 21508 15852 21514 15904
rect 22066 15892 22094 15932
rect 23750 15892 23756 15904
rect 22066 15864 23756 15892
rect 23750 15852 23756 15864
rect 23808 15852 23814 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 9088 15660 9137 15688
rect 9088 15648 9094 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 11609 15691 11667 15697
rect 11609 15657 11621 15691
rect 11655 15688 11667 15691
rect 11698 15688 11704 15700
rect 11655 15660 11704 15688
rect 11655 15657 11667 15660
rect 11609 15651 11667 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 14458 15688 14464 15700
rect 12676 15660 14464 15688
rect 12676 15648 12682 15660
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 16390 15648 16396 15700
rect 16448 15648 16454 15700
rect 17310 15688 17316 15700
rect 16868 15660 17316 15688
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 13446 15620 13452 15632
rect 12032 15592 13452 15620
rect 12032 15580 12038 15592
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 15010 15580 15016 15632
rect 15068 15620 15074 15632
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 15068 15592 15485 15620
rect 15068 15580 15074 15592
rect 15473 15589 15485 15592
rect 15519 15620 15531 15623
rect 16868 15620 16896 15660
rect 17310 15648 17316 15660
rect 17368 15688 17374 15700
rect 18506 15688 18512 15700
rect 17368 15660 18512 15688
rect 17368 15648 17374 15660
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 21450 15648 21456 15700
rect 21508 15688 21514 15700
rect 24946 15688 24952 15700
rect 21508 15660 24952 15688
rect 21508 15648 21514 15660
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 15519 15592 16896 15620
rect 21821 15623 21879 15629
rect 15519 15589 15531 15592
rect 15473 15583 15531 15589
rect 21821 15589 21833 15623
rect 21867 15620 21879 15623
rect 22738 15620 22744 15632
rect 21867 15592 22744 15620
rect 21867 15589 21879 15592
rect 21821 15583 21879 15589
rect 22738 15580 22744 15592
rect 22796 15580 22802 15632
rect 24118 15580 24124 15632
rect 24176 15620 24182 15632
rect 25041 15623 25099 15629
rect 25041 15620 25053 15623
rect 24176 15592 25053 15620
rect 24176 15580 24182 15592
rect 25041 15589 25053 15592
rect 25087 15620 25099 15623
rect 25225 15623 25283 15629
rect 25225 15620 25237 15623
rect 25087 15592 25237 15620
rect 25087 15589 25099 15592
rect 25041 15583 25099 15589
rect 25225 15589 25237 15592
rect 25271 15589 25283 15623
rect 25225 15583 25283 15589
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 6886 15524 9689 15552
rect 6886 15496 6914 15524
rect 9677 15521 9689 15524
rect 9723 15552 9735 15555
rect 10686 15552 10692 15564
rect 9723 15524 10692 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 11940 15524 12173 15552
rect 11940 15512 11946 15524
rect 12161 15521 12173 15524
rect 12207 15552 12219 15555
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12207 15524 12633 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18598 15552 18604 15564
rect 18187 15524 18604 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 20254 15552 20260 15564
rect 19475 15524 20260 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 20772 15524 21680 15552
rect 20772 15512 20778 15524
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 6822 15484 6828 15496
rect 6604 15456 6828 15484
rect 6604 15444 6610 15456
rect 6822 15444 6828 15456
rect 6880 15456 6914 15496
rect 6880 15444 6886 15456
rect 9490 15444 9496 15496
rect 9548 15484 9554 15496
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9548 15456 9597 15484
rect 9548 15444 9554 15456
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15484 10287 15487
rect 12250 15484 12256 15496
rect 10275 15456 12256 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 21652 15493 21680 15524
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22278 15552 22284 15564
rect 22152 15524 22284 15552
rect 22152 15512 22158 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 23658 15512 23664 15564
rect 23716 15552 23722 15564
rect 24029 15555 24087 15561
rect 24029 15552 24041 15555
rect 23716 15524 24041 15552
rect 23716 15512 23722 15524
rect 24029 15521 24041 15524
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 24762 15512 24768 15564
rect 24820 15512 24826 15564
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12618 15416 12624 15428
rect 12023 15388 12624 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 17865 15419 17923 15425
rect 17434 15388 17540 15416
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 9493 15351 9551 15357
rect 9493 15348 9505 15351
rect 9456 15320 9505 15348
rect 9456 15308 9462 15320
rect 9493 15317 9505 15320
rect 9539 15317 9551 15351
rect 9493 15311 9551 15317
rect 12066 15308 12072 15360
rect 12124 15308 12130 15360
rect 13265 15351 13323 15357
rect 13265 15317 13277 15351
rect 13311 15348 13323 15351
rect 13722 15348 13728 15360
rect 13311 15320 13728 15348
rect 13311 15317 13323 15320
rect 13265 15311 13323 15317
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 15930 15308 15936 15360
rect 15988 15308 15994 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 17512 15348 17540 15388
rect 17865 15385 17877 15419
rect 17911 15416 17923 15419
rect 18322 15416 18328 15428
rect 17911 15388 18328 15416
rect 17911 15385 17923 15388
rect 17865 15379 17923 15385
rect 18322 15376 18328 15388
rect 18380 15376 18386 15428
rect 19610 15376 19616 15428
rect 19668 15416 19674 15428
rect 19705 15419 19763 15425
rect 19705 15416 19717 15419
rect 19668 15388 19717 15416
rect 19668 15376 19674 15388
rect 19705 15385 19717 15388
rect 19751 15385 19763 15419
rect 21266 15416 21272 15428
rect 20930 15388 21272 15416
rect 19705 15379 19763 15385
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22244 15388 22586 15416
rect 22244 15376 22250 15388
rect 23750 15376 23756 15428
rect 23808 15376 23814 15428
rect 18509 15351 18567 15357
rect 18509 15348 18521 15351
rect 16908 15320 18521 15348
rect 16908 15308 16914 15320
rect 18509 15317 18521 15320
rect 18555 15348 18567 15351
rect 19058 15348 19064 15360
rect 18555 15320 19064 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20530 15348 20536 15360
rect 19852 15320 20536 15348
rect 19852 15308 19858 15320
rect 20530 15308 20536 15320
rect 20588 15348 20594 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 20588 15320 21189 15348
rect 20588 15308 20594 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10008 15116 10149 15144
rect 10008 15104 10014 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 11330 15104 11336 15156
rect 11388 15104 11394 15156
rect 12161 15147 12219 15153
rect 12161 15113 12173 15147
rect 12207 15144 12219 15147
rect 12250 15144 12256 15156
rect 12207 15116 12256 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14274 15144 14280 15156
rect 14139 15116 14280 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14461 15147 14519 15153
rect 14461 15113 14473 15147
rect 14507 15113 14519 15147
rect 14461 15107 14519 15113
rect 8662 15036 8668 15088
rect 8720 15036 8726 15088
rect 14476 15076 14504 15107
rect 15930 15104 15936 15156
rect 15988 15104 15994 15156
rect 16298 15104 16304 15156
rect 16356 15104 16362 15156
rect 17402 15104 17408 15156
rect 17460 15144 17466 15156
rect 17497 15147 17555 15153
rect 17497 15144 17509 15147
rect 17460 15116 17509 15144
rect 17460 15104 17466 15116
rect 17497 15113 17509 15116
rect 17543 15113 17555 15147
rect 17497 15107 17555 15113
rect 19886 15104 19892 15156
rect 19944 15104 19950 15156
rect 20809 15147 20867 15153
rect 20809 15113 20821 15147
rect 20855 15144 20867 15147
rect 21818 15144 21824 15156
rect 20855 15116 21824 15144
rect 20855 15113 20867 15116
rect 20809 15107 20867 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 17034 15076 17040 15088
rect 9692 15048 14412 15076
rect 14476 15048 17040 15076
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 6880 14912 7665 14940
rect 6880 14900 6886 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8294 14940 8300 14952
rect 7975 14912 8300 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 9692 14949 9720 15048
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 11606 15008 11612 15020
rect 10643 14980 11612 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13372 14980 14013 15008
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9364 14912 9689 14940
rect 9364 14900 9370 14912
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 10686 14900 10692 14952
rect 10744 14900 10750 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13372 14949 13400 14980
rect 14001 14977 14013 14980
rect 14047 14977 14059 15011
rect 14384 15008 14412 15048
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 18785 15079 18843 15085
rect 18785 15045 18797 15079
rect 18831 15076 18843 15079
rect 20070 15076 20076 15088
rect 18831 15048 20076 15076
rect 18831 15045 18843 15048
rect 18785 15039 18843 15045
rect 20070 15036 20076 15048
rect 20128 15036 20134 15088
rect 22830 15076 22836 15088
rect 21008 15048 22836 15076
rect 15194 15008 15200 15020
rect 14384 14980 15200 15008
rect 14001 14971 14059 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 16942 15008 16948 15020
rect 15764 14980 16948 15008
rect 13357 14943 13415 14949
rect 13357 14940 13369 14943
rect 12492 14912 13369 14940
rect 12492 14900 12498 14912
rect 13357 14909 13369 14912
rect 13403 14909 13415 14943
rect 13357 14903 13415 14909
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 14550 14940 14556 14952
rect 13955 14912 14556 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 15764 14949 15792 14980
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 18874 14968 18880 15020
rect 18932 15008 18938 15020
rect 21008 15017 21036 15048
rect 22830 15036 22836 15048
rect 22888 15036 22894 15088
rect 23290 15036 23296 15088
rect 23348 15036 23354 15088
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 18932 14980 19993 15008
rect 18932 14968 18938 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21266 14968 21272 15020
rect 21324 14968 21330 15020
rect 22094 14968 22100 15020
rect 22152 14968 22158 15020
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 15841 14943 15899 14949
rect 15841 14909 15853 14943
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 12526 14764 12532 14816
rect 12584 14764 12590 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15470 14804 15476 14816
rect 15335 14776 15476 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15470 14764 15476 14776
rect 15528 14804 15534 14816
rect 15856 14804 15884 14903
rect 19794 14900 19800 14952
rect 19852 14900 19858 14952
rect 21284 14940 21312 14968
rect 20272 14912 21312 14940
rect 18598 14832 18604 14884
rect 18656 14832 18662 14884
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 20272 14872 20300 14912
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 19116 14844 20300 14872
rect 20349 14875 20407 14881
rect 19116 14832 19122 14844
rect 20349 14841 20361 14875
rect 20395 14872 20407 14875
rect 22830 14872 22836 14884
rect 20395 14844 22836 14872
rect 20395 14841 20407 14844
rect 20349 14835 20407 14841
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 15528 14776 15884 14804
rect 15528 14764 15534 14776
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7892 14572 8217 14600
rect 7892 14560 7898 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13173 14603 13231 14609
rect 13173 14600 13185 14603
rect 12860 14572 13185 14600
rect 12860 14560 12866 14572
rect 13173 14569 13185 14572
rect 13219 14569 13231 14603
rect 13173 14563 13231 14569
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 24302 14600 24308 14612
rect 20772 14572 24308 14600
rect 20772 14560 20778 14572
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 15378 14492 15384 14544
rect 15436 14532 15442 14544
rect 20806 14532 20812 14544
rect 15436 14504 20812 14532
rect 15436 14492 15442 14504
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 22002 14532 22008 14544
rect 21192 14504 22008 14532
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 7282 14464 7288 14476
rect 6779 14436 7288 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 6472 14328 6500 14427
rect 7282 14424 7288 14436
rect 7340 14424 7346 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11296 14436 11989 14464
rect 11296 14424 11302 14436
rect 11977 14433 11989 14436
rect 12023 14464 12035 14467
rect 12250 14464 12256 14476
rect 12023 14436 12256 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12250 14424 12256 14436
rect 12308 14464 12314 14476
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12308 14436 12541 14464
rect 12308 14424 12314 14436
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 12529 14427 12587 14433
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 13044 14436 13553 14464
rect 13044 14424 13050 14436
rect 13541 14433 13553 14436
rect 13587 14464 13599 14467
rect 14921 14467 14979 14473
rect 13587 14436 14872 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9640 14368 9965 14396
rect 9640 14356 9646 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14734 14396 14740 14408
rect 13872 14368 14740 14396
rect 13872 14356 13878 14368
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 14844 14396 14872 14436
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15194 14464 15200 14476
rect 14967 14436 15200 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 16022 14424 16028 14476
rect 16080 14464 16086 14476
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16080 14436 16589 14464
rect 16080 14424 16086 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 19886 14396 19892 14408
rect 14844 14368 19892 14396
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14392 20499 14399
rect 21192 14396 21220 14504
rect 22002 14492 22008 14504
rect 22060 14492 22066 14544
rect 23934 14492 23940 14544
rect 23992 14532 23998 14544
rect 23992 14504 25084 14532
rect 23992 14492 23998 14504
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14433 21695 14467
rect 21637 14427 21695 14433
rect 20548 14392 21220 14396
rect 20487 14368 21220 14392
rect 21652 14396 21680 14427
rect 21726 14424 21732 14476
rect 21784 14424 21790 14476
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 24854 14464 24860 14476
rect 23431 14436 24860 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 23290 14396 23296 14408
rect 21652 14368 23296 14396
rect 20487 14365 20576 14368
rect 20441 14364 20576 14365
rect 20441 14359 20499 14364
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 24029 14399 24087 14405
rect 24029 14365 24041 14399
rect 24075 14396 24087 14399
rect 24486 14396 24492 14408
rect 24075 14368 24492 14396
rect 24075 14365 24087 14368
rect 24029 14359 24087 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 25056 14405 25084 14504
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14365 25099 14399
rect 25041 14359 25099 14365
rect 6822 14328 6828 14340
rect 6472 14300 6828 14328
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 7958 14300 8616 14328
rect 8588 14269 8616 14300
rect 10134 14288 10140 14340
rect 10192 14328 10198 14340
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 10192 14300 10241 14328
rect 10192 14288 10198 14300
rect 10229 14297 10241 14300
rect 10275 14297 10287 14331
rect 12158 14328 12164 14340
rect 11454 14300 12164 14328
rect 10229 14291 10287 14297
rect 8573 14263 8631 14269
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 8662 14260 8668 14272
rect 8619 14232 8668 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9677 14263 9735 14269
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 11238 14260 11244 14272
rect 9723 14232 11244 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 11238 14220 11244 14232
rect 11296 14260 11302 14272
rect 11532 14260 11560 14300
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 12713 14331 12771 14337
rect 12713 14297 12725 14331
rect 12759 14328 12771 14331
rect 14182 14328 14188 14340
rect 12759 14300 14188 14328
rect 12759 14297 12771 14300
rect 12713 14291 12771 14297
rect 14182 14288 14188 14300
rect 14240 14288 14246 14340
rect 14645 14331 14703 14337
rect 14645 14297 14657 14331
rect 14691 14328 14703 14331
rect 15378 14328 15384 14340
rect 14691 14300 15384 14328
rect 14691 14297 14703 14300
rect 14645 14291 14703 14297
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 16853 14331 16911 14337
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 16899 14300 17693 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17681 14297 17693 14300
rect 17727 14297 17739 14331
rect 17681 14291 17739 14297
rect 19610 14288 19616 14340
rect 19668 14328 19674 14340
rect 23382 14328 23388 14340
rect 19668 14300 23388 14328
rect 19668 14288 19674 14300
rect 23382 14288 23388 14300
rect 23440 14288 23446 14340
rect 11296 14232 11560 14260
rect 11296 14220 11302 14232
rect 12802 14220 12808 14272
rect 12860 14220 12866 14272
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 14366 14260 14372 14272
rect 14323 14232 14372 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 16761 14263 16819 14269
rect 16761 14260 16773 14263
rect 15712 14232 16773 14260
rect 15712 14220 15718 14232
rect 16761 14229 16773 14232
rect 16807 14229 16819 14263
rect 16761 14223 16819 14229
rect 17221 14263 17279 14269
rect 17221 14229 17233 14263
rect 17267 14260 17279 14263
rect 20162 14260 20168 14272
rect 17267 14232 20168 14260
rect 17267 14229 17279 14232
rect 17221 14223 17279 14229
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 20254 14220 20260 14272
rect 20312 14220 20318 14272
rect 20438 14220 20444 14272
rect 20496 14260 20502 14272
rect 21821 14263 21879 14269
rect 21821 14260 21833 14263
rect 20496 14232 21833 14260
rect 20496 14220 20502 14232
rect 21821 14229 21833 14232
rect 21867 14229 21879 14263
rect 21821 14223 21879 14229
rect 22189 14263 22247 14269
rect 22189 14229 22201 14263
rect 22235 14260 22247 14263
rect 23934 14260 23940 14272
rect 22235 14232 23940 14260
rect 22235 14229 22247 14232
rect 22189 14223 22247 14229
rect 23934 14220 23940 14232
rect 23992 14220 23998 14272
rect 24857 14263 24915 14269
rect 24857 14229 24869 14263
rect 24903 14260 24915 14263
rect 25130 14260 25136 14272
rect 24903 14232 25136 14260
rect 24903 14229 24915 14232
rect 24857 14223 24915 14229
rect 25130 14220 25136 14232
rect 25188 14220 25194 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 9916 14028 12633 14056
rect 9916 14016 9922 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 12986 14016 12992 14068
rect 13044 14016 13050 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 15565 14059 15623 14065
rect 14792 14028 15424 14056
rect 14792 14016 14798 14028
rect 8294 13988 8300 14000
rect 7760 13960 8300 13988
rect 6822 13880 6828 13932
rect 6880 13920 6886 13932
rect 7760 13929 7788 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8662 13948 8668 14000
rect 8720 13948 8726 14000
rect 11149 13991 11207 13997
rect 11149 13957 11161 13991
rect 11195 13988 11207 13991
rect 11330 13988 11336 14000
rect 11195 13960 11336 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 11330 13948 11336 13960
rect 11388 13948 11394 14000
rect 12250 13948 12256 14000
rect 12308 13948 12314 14000
rect 15396 13988 15424 14028
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16022 14056 16028 14068
rect 15611 14028 16028 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 18601 14059 18659 14065
rect 16132 14028 18460 14056
rect 16132 13988 16160 14028
rect 15396 13960 16160 13988
rect 18432 13988 18460 14028
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18782 14056 18788 14068
rect 18647 14028 18788 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19058 14016 19064 14068
rect 19116 14016 19122 14068
rect 20349 14059 20407 14065
rect 20349 14025 20361 14059
rect 20395 14056 20407 14059
rect 21174 14056 21180 14068
rect 20395 14028 21180 14056
rect 20395 14025 20407 14028
rect 20349 14019 20407 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 22189 14059 22247 14065
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 22646 14056 22652 14068
rect 22235 14028 22652 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 24084 14028 25053 14056
rect 24084 14016 24090 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 18432 13960 19441 13988
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 19610 13948 19616 14000
rect 19668 13948 19674 14000
rect 22462 13988 22468 14000
rect 21100 13960 22468 13988
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 6880 13892 7757 13920
rect 6880 13880 6886 13892
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 9582 13920 9588 13932
rect 7745 13883 7803 13889
rect 9232 13892 9588 13920
rect 8018 13812 8024 13864
rect 8076 13812 8082 13864
rect 9030 13812 9036 13864
rect 9088 13852 9094 13864
rect 9232 13852 9260 13892
rect 9582 13880 9588 13892
rect 9640 13920 9646 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 9640 13892 10333 13920
rect 9640 13880 9646 13892
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 11882 13920 11888 13932
rect 10321 13883 10379 13889
rect 11624 13892 11888 13920
rect 9088 13824 9260 13852
rect 9769 13855 9827 13861
rect 9088 13812 9094 13824
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10134 13852 10140 13864
rect 9815 13824 10140 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10134 13812 10140 13824
rect 10192 13852 10198 13864
rect 11624 13852 11652 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 19058 13920 19064 13932
rect 12584 13892 13216 13920
rect 15226 13892 15976 13920
rect 12584 13880 12590 13892
rect 10192 13824 11652 13852
rect 10192 13812 10198 13824
rect 11698 13812 11704 13864
rect 11756 13812 11762 13864
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13188 13861 13216 13892
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12768 13824 13093 13852
rect 12768 13812 12774 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 13188 13784 13216 13815
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 15948 13861 15976 13892
rect 18156 13892 19064 13920
rect 15933 13855 15991 13861
rect 13924 13824 15148 13852
rect 13924 13784 13952 13824
rect 13188 13756 13952 13784
rect 15120 13784 15148 13824
rect 15933 13821 15945 13855
rect 15979 13852 15991 13855
rect 16482 13852 16488 13864
rect 15979 13824 16488 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 16482 13812 16488 13824
rect 16540 13852 16546 13864
rect 16540 13824 16804 13852
rect 16540 13812 16546 13824
rect 15194 13784 15200 13796
rect 15120 13756 15200 13784
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 16776 13784 16804 13824
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 18156 13852 18184 13892
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 20162 13880 20168 13932
rect 20220 13880 20226 13932
rect 21100 13929 21128 13960
rect 22462 13948 22468 13960
rect 22520 13948 22526 14000
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 22002 13880 22008 13932
rect 22060 13880 22066 13932
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 25225 13923 25283 13929
rect 25225 13920 25237 13923
rect 24452 13892 25237 13920
rect 24452 13880 24458 13892
rect 25225 13889 25237 13892
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 16960 13824 18184 13852
rect 18248 13824 18889 13852
rect 16960 13784 16988 13824
rect 18248 13784 18276 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 21266 13852 21272 13864
rect 18877 13815 18935 13821
rect 20916 13824 21272 13852
rect 16776 13756 16988 13784
rect 18156 13756 18276 13784
rect 14090 13725 14096 13728
rect 14080 13719 14096 13725
rect 14080 13685 14092 13719
rect 14080 13679 14096 13685
rect 14090 13676 14096 13679
rect 14148 13676 14154 13728
rect 17116 13719 17174 13725
rect 17116 13685 17128 13719
rect 17162 13716 17174 13719
rect 17310 13716 17316 13728
rect 17162 13688 17316 13716
rect 17162 13685 17174 13688
rect 17116 13679 17174 13685
rect 17310 13676 17316 13688
rect 17368 13716 17374 13728
rect 17586 13716 17592 13728
rect 17368 13688 17592 13716
rect 17368 13676 17374 13688
rect 17586 13676 17592 13688
rect 17644 13716 17650 13728
rect 18156 13716 18184 13756
rect 18506 13744 18512 13796
rect 18564 13784 18570 13796
rect 20916 13793 20944 13824
rect 21266 13812 21272 13824
rect 21324 13812 21330 13864
rect 22186 13812 22192 13864
rect 22244 13852 22250 13864
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22244 13824 22845 13852
rect 22244 13812 22250 13824
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 23198 13812 23204 13864
rect 23256 13852 23262 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 23256 13824 24593 13852
rect 23256 13812 23262 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 20901 13787 20959 13793
rect 18564 13756 19196 13784
rect 18564 13744 18570 13756
rect 17644 13688 18184 13716
rect 19168 13716 19196 13756
rect 20901 13753 20913 13787
rect 20947 13753 20959 13787
rect 20901 13747 20959 13753
rect 20990 13716 20996 13728
rect 19168 13688 20996 13716
rect 17644 13676 17650 13688
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 22278 13676 22284 13728
rect 22336 13716 22342 13728
rect 22646 13716 22652 13728
rect 22336 13688 22652 13716
rect 22336 13676 22342 13688
rect 22646 13676 22652 13688
rect 22704 13716 22710 13728
rect 23090 13719 23148 13725
rect 23090 13716 23102 13719
rect 22704 13688 23102 13716
rect 22704 13676 22710 13688
rect 23090 13685 23102 13688
rect 23136 13685 23148 13719
rect 23090 13679 23148 13685
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 6546 13472 6552 13524
rect 6604 13472 6610 13524
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 7708 13484 9229 13512
rect 7708 13472 7714 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 13906 13472 13912 13524
rect 13964 13472 13970 13524
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 15654 13512 15660 13524
rect 14608 13484 15660 13512
rect 14608 13472 14614 13484
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 15746 13472 15752 13524
rect 15804 13472 15810 13524
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 17402 13512 17408 13524
rect 16724 13484 17408 13512
rect 16724 13472 16730 13484
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 24210 13512 24216 13524
rect 17644 13484 24216 13512
rect 17644 13472 17650 13484
rect 24210 13472 24216 13484
rect 24268 13472 24274 13524
rect 24486 13472 24492 13524
rect 24544 13512 24550 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24544 13484 24593 13512
rect 24544 13472 24550 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 15562 13444 15568 13456
rect 13320 13416 15568 13444
rect 13320 13404 13326 13416
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 15764 13444 15792 13472
rect 21082 13444 21088 13456
rect 15764 13416 21088 13444
rect 21082 13404 21088 13416
rect 21140 13404 21146 13456
rect 21174 13404 21180 13456
rect 21232 13444 21238 13456
rect 21232 13416 24808 13444
rect 21232 13404 21238 13416
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 7340 13348 9781 13376
rect 7340 13336 7346 13348
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 12161 13379 12219 13385
rect 12161 13376 12173 13379
rect 11572 13348 12173 13376
rect 11572 13336 11578 13348
rect 12161 13345 12173 13348
rect 12207 13376 12219 13379
rect 13449 13379 13507 13385
rect 13449 13376 13461 13379
rect 12207 13348 13461 13376
rect 12207 13345 12219 13348
rect 12161 13339 12219 13345
rect 13449 13345 13461 13348
rect 13495 13376 13507 13379
rect 13814 13376 13820 13388
rect 13495 13348 13820 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15344 13348 15761 13376
rect 15344 13336 15350 13348
rect 15749 13345 15761 13348
rect 15795 13376 15807 13379
rect 15930 13376 15936 13388
rect 15795 13348 15936 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 20070 13376 20076 13388
rect 16347 13348 20076 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 9030 13308 9036 13320
rect 8352 13280 9036 13308
rect 8352 13268 8358 13280
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13308 12679 13311
rect 13906 13308 13912 13320
rect 12667 13280 13912 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 14976 13280 15669 13308
rect 14976 13268 14982 13280
rect 15657 13277 15669 13280
rect 15703 13308 15715 13311
rect 16114 13308 16120 13320
rect 15703 13280 16120 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 8021 13243 8079 13249
rect 7590 13212 7972 13240
rect 7944 13172 7972 13212
rect 8021 13209 8033 13243
rect 8067 13240 8079 13243
rect 9122 13240 9128 13252
rect 8067 13212 9128 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 9631 13212 10640 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 8662 13172 8668 13184
rect 7944 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 10612 13172 10640 13212
rect 11238 13200 11244 13252
rect 11296 13200 11302 13252
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 11885 13243 11943 13249
rect 11885 13240 11897 13243
rect 11848 13212 11897 13240
rect 11848 13200 11854 13212
rect 11885 13209 11897 13212
rect 11931 13209 11943 13243
rect 11885 13203 11943 13209
rect 12158 13200 12164 13252
rect 12216 13240 12222 13252
rect 14645 13243 14703 13249
rect 14645 13240 14657 13243
rect 12216 13212 14657 13240
rect 12216 13200 12222 13212
rect 14645 13209 14657 13212
rect 14691 13240 14703 13243
rect 15470 13240 15476 13252
rect 14691 13212 15476 13240
rect 14691 13209 14703 13212
rect 14645 13203 14703 13209
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 15565 13243 15623 13249
rect 15565 13209 15577 13243
rect 15611 13240 15623 13243
rect 16316 13240 16344 13339
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 23382 13336 23388 13388
rect 23440 13336 23446 13388
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17460 13280 17969 13308
rect 17460 13268 17466 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18693 13311 18751 13317
rect 18693 13308 18705 13311
rect 18380 13280 18705 13308
rect 18380 13268 18386 13280
rect 18693 13277 18705 13280
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 15611 13212 16344 13240
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17773 13243 17831 13249
rect 17773 13240 17785 13243
rect 17092 13212 17785 13240
rect 17092 13200 17098 13212
rect 17773 13209 17785 13212
rect 17819 13209 17831 13243
rect 17773 13203 17831 13209
rect 18506 13200 18512 13252
rect 18564 13200 18570 13252
rect 12342 13172 12348 13184
rect 10612 13144 12348 13172
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 14918 13132 14924 13184
rect 14976 13132 14982 13184
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 18708 13172 18736 13271
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19392 13280 19441 13308
rect 19392 13268 19398 13280
rect 19429 13277 19441 13280
rect 19475 13308 19487 13311
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 19475 13280 20821 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21910 13268 21916 13320
rect 21968 13268 21974 13320
rect 22189 13311 22247 13317
rect 22189 13277 22201 13311
rect 22235 13277 22247 13311
rect 22189 13271 22247 13277
rect 20257 13243 20315 13249
rect 20257 13209 20269 13243
rect 20303 13240 20315 13243
rect 22204 13240 22232 13271
rect 24026 13268 24032 13320
rect 24084 13268 24090 13320
rect 24780 13317 24808 13416
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 24302 13240 24308 13252
rect 20303 13212 22094 13240
rect 22204 13212 24308 13240
rect 20303 13209 20315 13212
rect 20257 13203 20315 13209
rect 20714 13172 20720 13184
rect 18708 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22066 13172 22094 13212
rect 24302 13200 24308 13212
rect 24360 13200 24366 13252
rect 24394 13200 24400 13252
rect 24452 13240 24458 13252
rect 25041 13243 25099 13249
rect 25041 13240 25053 13243
rect 24452 13212 25053 13240
rect 24452 13200 24458 13212
rect 25041 13209 25053 13212
rect 25087 13209 25099 13243
rect 25041 13203 25099 13209
rect 22186 13172 22192 13184
rect 22066 13144 22192 13172
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 7377 12971 7435 12977
rect 7377 12937 7389 12971
rect 7423 12968 7435 12971
rect 7558 12968 7564 12980
rect 7423 12940 7564 12968
rect 7423 12937 7435 12940
rect 7377 12931 7435 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 9490 12928 9496 12980
rect 9548 12968 9554 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9548 12940 9781 12968
rect 9548 12928 9554 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 9769 12931 9827 12937
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 11698 12968 11704 12980
rect 10827 12940 11704 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12250 12968 12256 12980
rect 12023 12940 12256 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 13354 12928 13360 12980
rect 13412 12928 13418 12980
rect 14550 12928 14556 12980
rect 14608 12928 14614 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14884 12940 15025 12968
rect 14884 12928 14890 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 17126 12928 17132 12980
rect 17184 12928 17190 12980
rect 17586 12928 17592 12980
rect 17644 12928 17650 12980
rect 18233 12971 18291 12977
rect 18233 12937 18245 12971
rect 18279 12937 18291 12971
rect 18233 12931 18291 12937
rect 6914 12900 6920 12912
rect 6886 12860 6920 12900
rect 6972 12860 6978 12912
rect 9309 12903 9367 12909
rect 9309 12869 9321 12903
rect 9355 12900 9367 12903
rect 9858 12900 9864 12912
rect 9355 12872 9864 12900
rect 9355 12869 9367 12872
rect 9309 12863 9367 12869
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 10873 12903 10931 12909
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 10919 12872 11192 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 6886 12832 6914 12860
rect 6840 12804 6914 12832
rect 7009 12835 7067 12841
rect 6840 12773 6868 12804
rect 7009 12801 7021 12835
rect 7055 12832 7067 12835
rect 7374 12832 7380 12844
rect 7055 12804 7380 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 7892 12804 8125 12832
rect 7892 12792 7898 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8996 12804 9413 12832
rect 8996 12792 9002 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 11164 12832 11192 12872
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 11296 12872 12081 12900
rect 11296 12860 11302 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 12069 12863 12127 12869
rect 12989 12903 13047 12909
rect 12989 12869 13001 12903
rect 13035 12900 13047 12903
rect 15562 12900 15568 12912
rect 13035 12872 14964 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 9401 12795 9459 12801
rect 10796 12804 11008 12832
rect 11164 12804 11621 12832
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12764 6975 12767
rect 8021 12767 8079 12773
rect 6963 12736 7052 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 7024 12708 7052 12736
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8478 12764 8484 12776
rect 8067 12736 8484 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 10042 12764 10048 12776
rect 9180 12736 10048 12764
rect 9180 12724 9186 12736
rect 10042 12724 10048 12736
rect 10100 12764 10106 12776
rect 10796 12764 10824 12804
rect 10980 12776 11008 12804
rect 11609 12801 11621 12804
rect 11655 12832 11667 12835
rect 13262 12832 13268 12844
rect 11655 12804 13268 12832
rect 11655 12801 11667 12804
rect 11609 12795 11667 12801
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13688 12804 14197 12832
rect 13688 12792 13694 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14936 12832 14964 12872
rect 15304 12872 15568 12900
rect 15304 12832 15332 12872
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 18248 12900 18276 12931
rect 19058 12928 19064 12980
rect 19116 12928 19122 12980
rect 19521 12971 19579 12977
rect 19521 12937 19533 12971
rect 19567 12968 19579 12971
rect 19978 12968 19984 12980
rect 19567 12940 19984 12968
rect 19567 12937 19579 12940
rect 19521 12931 19579 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 22002 12968 22008 12980
rect 20088 12940 22008 12968
rect 20088 12900 20116 12940
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22189 12971 22247 12977
rect 22189 12968 22201 12971
rect 22152 12940 22201 12968
rect 22152 12928 22158 12940
rect 22189 12937 22201 12940
rect 22235 12937 22247 12971
rect 22189 12931 22247 12937
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 23474 12968 23480 12980
rect 22787 12940 23480 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 23474 12928 23480 12940
rect 23532 12968 23538 12980
rect 24394 12968 24400 12980
rect 23532 12940 24400 12968
rect 23532 12928 23538 12940
rect 22370 12900 22376 12912
rect 18248 12872 20116 12900
rect 20180 12872 22376 12900
rect 14936 12804 15332 12832
rect 15381 12835 15439 12841
rect 14185 12795 14243 12801
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 15427 12804 16160 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 10100 12736 10824 12764
rect 10100 12724 10106 12736
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 12250 12724 12256 12776
rect 12308 12764 12314 12776
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 12308 12736 12725 12764
rect 12308 12724 12314 12736
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 7006 12656 7012 12708
rect 7064 12656 7070 12708
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 9456 12668 10425 12696
rect 9456 12656 9462 12668
rect 10413 12665 10425 12668
rect 10459 12665 10471 12699
rect 10413 12659 10471 12665
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 11701 12699 11759 12705
rect 11701 12696 11713 12699
rect 10836 12668 11713 12696
rect 10836 12656 10842 12668
rect 11701 12665 11713 12668
rect 11747 12696 11759 12699
rect 12526 12696 12532 12708
rect 11747 12668 12532 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12912 12696 12940 12727
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 13998 12764 14004 12776
rect 13872 12736 14004 12764
rect 13872 12724 13878 12736
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 14093 12767 14151 12773
rect 14093 12733 14105 12767
rect 14139 12764 14151 12767
rect 15286 12764 15292 12776
rect 14139 12736 15292 12764
rect 14139 12733 14151 12736
rect 14093 12727 14151 12733
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 15528 12736 15577 12764
rect 15528 12724 15534 12736
rect 15565 12733 15577 12736
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 15378 12696 15384 12708
rect 12912 12668 15384 12696
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 16132 12705 16160 12804
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18322 12832 18328 12844
rect 18095 12804 18328 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 20180 12841 20208 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 23290 12860 23296 12912
rect 23348 12900 23354 12912
rect 23385 12903 23443 12909
rect 23385 12900 23397 12903
rect 23348 12872 23397 12900
rect 23348 12860 23354 12872
rect 23385 12869 23397 12872
rect 23431 12869 23443 12903
rect 23768 12900 23796 12940
rect 24394 12928 24400 12940
rect 24452 12968 24458 12980
rect 25133 12971 25191 12977
rect 25133 12968 25145 12971
rect 24452 12940 25145 12968
rect 24452 12928 24458 12940
rect 25133 12937 25145 12940
rect 25179 12937 25191 12971
rect 25133 12931 25191 12937
rect 23768 12872 23874 12900
rect 23385 12863 23443 12869
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 20622 12792 20628 12844
rect 20680 12792 20686 12844
rect 21082 12792 21088 12844
rect 21140 12792 21146 12844
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12832 22063 12835
rect 22094 12832 22100 12844
rect 22051 12804 22100 12832
rect 22051 12801 22063 12804
rect 22005 12795 22063 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22244 12804 23121 12832
rect 22244 12792 22250 12804
rect 23109 12801 23121 12804
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12764 17095 12767
rect 18782 12764 18788 12776
rect 17083 12736 18788 12764
rect 17083 12733 17095 12736
rect 17037 12727 17095 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 18969 12767 19027 12773
rect 18969 12733 18981 12767
rect 19015 12764 19027 12767
rect 20640 12764 20668 12792
rect 19015 12736 20668 12764
rect 20901 12767 20959 12773
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 20901 12733 20913 12767
rect 20947 12733 20959 12767
rect 20901 12727 20959 12733
rect 16117 12699 16175 12705
rect 16117 12665 16129 12699
rect 16163 12696 16175 12699
rect 20622 12696 20628 12708
rect 16163 12668 20628 12696
rect 16163 12665 16175 12668
rect 16117 12659 16175 12665
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 20916 12696 20944 12727
rect 20990 12724 20996 12776
rect 21048 12764 21054 12776
rect 22465 12767 22523 12773
rect 22465 12764 22477 12767
rect 21048 12736 22477 12764
rect 21048 12724 21054 12736
rect 22465 12733 22477 12736
rect 22511 12733 22523 12767
rect 22465 12727 22523 12733
rect 20916 12668 23244 12696
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12628 8631 12631
rect 11146 12628 11152 12640
rect 8619 12600 11152 12628
rect 8619 12597 8631 12600
rect 8573 12591 8631 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11848 12600 12265 12628
rect 11848 12588 11854 12600
rect 12253 12597 12265 12600
rect 12299 12628 12311 12631
rect 12710 12628 12716 12640
rect 12299 12600 12716 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 13504 12600 19993 12628
rect 13504 12588 13510 12600
rect 19981 12597 19993 12600
rect 20027 12597 20039 12631
rect 19981 12591 20039 12597
rect 21450 12588 21456 12640
rect 21508 12588 21514 12640
rect 23216 12628 23244 12668
rect 23382 12628 23388 12640
rect 23216 12600 23388 12628
rect 23382 12588 23388 12600
rect 23440 12628 23446 12640
rect 24857 12631 24915 12637
rect 24857 12628 24869 12631
rect 23440 12600 24869 12628
rect 23440 12588 23446 12600
rect 24857 12597 24869 12600
rect 24903 12597 24915 12631
rect 24857 12591 24915 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 10226 12384 10232 12436
rect 10284 12384 10290 12436
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 10560 12396 11437 12424
rect 10560 12384 10566 12396
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12032 12396 12572 12424
rect 12032 12384 12038 12396
rect 12434 12356 12440 12368
rect 10704 12328 12440 12356
rect 7374 12248 7380 12300
rect 7432 12248 7438 12300
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 10704 12297 10732 12328
rect 12434 12316 12440 12328
rect 12492 12316 12498 12368
rect 12544 12356 12572 12396
rect 12618 12384 12624 12436
rect 12676 12384 12682 12436
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 13596 12396 13768 12424
rect 13596 12384 13602 12396
rect 12710 12356 12716 12368
rect 12544 12328 12716 12356
rect 12710 12316 12716 12328
rect 12768 12316 12774 12368
rect 13633 12359 13691 12365
rect 13633 12356 13645 12359
rect 13096 12328 13645 12356
rect 13096 12300 13124 12328
rect 13633 12325 13645 12328
rect 13679 12325 13691 12359
rect 13633 12319 13691 12325
rect 13740 12356 13768 12396
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 14148 12396 14289 12424
rect 14148 12384 14154 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 14884 12396 14964 12424
rect 14884 12384 14890 12396
rect 13740 12328 14872 12356
rect 10689 12291 10747 12297
rect 10689 12257 10701 12291
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 10796 12220 10824 12251
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11020 12260 12081 12288
rect 11020 12248 11026 12260
rect 12069 12257 12081 12260
rect 12115 12288 12127 12291
rect 12158 12288 12164 12300
rect 12115 12260 12164 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 13078 12288 13084 12300
rect 12584 12260 13084 12288
rect 12584 12248 12590 12260
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13740 12288 13768 12328
rect 14844 12300 14872 12328
rect 13311 12260 13768 12288
rect 13909 12291 13967 12297
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13909 12257 13921 12291
rect 13955 12288 13967 12291
rect 13998 12288 14004 12300
rect 13955 12260 14004 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 13998 12248 14004 12260
rect 14056 12288 14062 12300
rect 14734 12288 14740 12300
rect 14056 12260 14740 12288
rect 14056 12248 14062 12260
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 14826 12248 14832 12300
rect 14884 12248 14890 12300
rect 7340 12192 10824 12220
rect 11793 12223 11851 12229
rect 7340 12180 7346 12192
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 14936 12220 14964 12396
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 18782 12424 18788 12436
rect 15344 12396 18788 12424
rect 15344 12384 15350 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19886 12424 19892 12436
rect 19484 12396 19892 12424
rect 19484 12384 19490 12396
rect 19886 12384 19892 12396
rect 19944 12424 19950 12436
rect 21358 12424 21364 12436
rect 19944 12396 21364 12424
rect 19944 12384 19950 12396
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24176 12396 24593 12424
rect 24176 12384 24182 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 15102 12316 15108 12368
rect 15160 12356 15166 12368
rect 15470 12356 15476 12368
rect 15160 12328 15476 12356
rect 15160 12316 15166 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 16022 12316 16028 12368
rect 16080 12356 16086 12368
rect 19058 12356 19064 12368
rect 16080 12328 19064 12356
rect 16080 12316 16086 12328
rect 19058 12316 19064 12328
rect 19116 12356 19122 12368
rect 19981 12359 20039 12365
rect 19981 12356 19993 12359
rect 19116 12328 19993 12356
rect 19116 12316 19122 12328
rect 19981 12325 19993 12328
rect 20027 12325 20039 12359
rect 19981 12319 20039 12325
rect 20254 12316 20260 12368
rect 20312 12356 20318 12368
rect 20530 12356 20536 12368
rect 20312 12328 20536 12356
rect 20312 12316 20318 12328
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 22554 12316 22560 12368
rect 22612 12356 22618 12368
rect 22830 12356 22836 12368
rect 22612 12328 22836 12356
rect 22612 12316 22618 12328
rect 22830 12316 22836 12328
rect 22888 12316 22894 12368
rect 18690 12288 18696 12300
rect 11839 12192 14964 12220
rect 15120 12260 18696 12288
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 10597 12155 10655 12161
rect 10597 12121 10609 12155
rect 10643 12152 10655 12155
rect 12526 12152 12532 12164
rect 10643 12124 12532 12152
rect 10643 12121 10655 12124
rect 10597 12115 10655 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 15120 12152 15148 12260
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 18877 12291 18935 12297
rect 18877 12257 18889 12291
rect 18923 12288 18935 12291
rect 19150 12288 19156 12300
rect 18923 12260 19156 12288
rect 18923 12257 18935 12260
rect 18877 12251 18935 12257
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 20714 12288 20720 12300
rect 19536 12260 20720 12288
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 16439 12192 18245 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 18233 12189 18245 12192
rect 18279 12220 18291 12223
rect 19334 12220 19340 12232
rect 18279 12192 19340 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 19536 12229 19564 12260
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 21266 12248 21272 12300
rect 21324 12288 21330 12300
rect 21913 12291 21971 12297
rect 21913 12288 21925 12291
rect 21324 12260 21925 12288
rect 21324 12248 21330 12260
rect 21913 12257 21925 12260
rect 21959 12257 21971 12291
rect 21913 12251 21971 12257
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12288 23443 12291
rect 24854 12288 24860 12300
rect 23431 12260 24860 12288
rect 23431 12257 23443 12260
rect 23385 12251 23443 12257
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22830 12220 22836 12232
rect 22244 12192 22836 12220
rect 22244 12180 22250 12192
rect 22830 12180 22836 12192
rect 22888 12180 22894 12232
rect 24026 12180 24032 12232
rect 24084 12180 24090 12232
rect 24118 12180 24124 12232
rect 24176 12220 24182 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24176 12192 24777 12220
rect 24176 12180 24182 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 14568 12124 15148 12152
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12710 12084 12716 12096
rect 11931 12056 12716 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13906 12084 13912 12096
rect 13035 12056 13912 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13906 12044 13912 12056
rect 13964 12084 13970 12096
rect 14568 12084 14596 12124
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17402 12152 17408 12164
rect 17000 12124 17408 12152
rect 17000 12112 17006 12124
rect 17402 12112 17408 12124
rect 17460 12112 17466 12164
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12152 19763 12155
rect 19886 12152 19892 12164
rect 19751 12124 19892 12152
rect 19751 12121 19763 12124
rect 19705 12115 19763 12121
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 21358 12112 21364 12164
rect 21416 12112 21422 12164
rect 13964 12056 14596 12084
rect 14645 12087 14703 12093
rect 13964 12044 13970 12056
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15378 12084 15384 12096
rect 14691 12056 15384 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15378 12044 15384 12056
rect 15436 12084 15442 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15436 12056 15669 12084
rect 15436 12044 15442 12056
rect 15657 12053 15669 12056
rect 15703 12084 15715 12087
rect 15838 12084 15844 12096
rect 15703 12056 15844 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 18414 12084 18420 12096
rect 16899 12056 18420 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 20346 12044 20352 12096
rect 20404 12084 20410 12096
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 20404 12056 20453 12084
rect 20404 12044 20410 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 7282 11840 7288 11892
rect 7340 11840 7346 11892
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 9582 11880 9588 11892
rect 8720 11852 9588 11880
rect 8720 11840 8726 11852
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9732 11852 9873 11880
rect 9732 11840 9738 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 11330 11880 11336 11892
rect 10284 11852 11336 11880
rect 10284 11840 10290 11852
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 12032 11852 12173 11880
rect 12032 11840 12038 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12161 11843 12219 11849
rect 12621 11883 12679 11889
rect 12621 11849 12633 11883
rect 12667 11880 12679 11883
rect 12802 11880 12808 11892
rect 12667 11852 12808 11880
rect 12667 11849 12679 11852
rect 12621 11843 12679 11849
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13078 11840 13084 11892
rect 13136 11880 13142 11892
rect 13538 11880 13544 11892
rect 13136 11852 13544 11880
rect 13136 11840 13142 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14458 11880 14464 11892
rect 14323 11852 14464 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 15654 11880 15660 11892
rect 14792 11852 15660 11880
rect 14792 11840 14798 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 17129 11883 17187 11889
rect 17129 11849 17141 11883
rect 17175 11880 17187 11883
rect 17494 11880 17500 11892
rect 17175 11852 17500 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 18325 11883 18383 11889
rect 18325 11880 18337 11883
rect 17920 11852 18337 11880
rect 17920 11840 17926 11852
rect 18325 11849 18337 11852
rect 18371 11849 18383 11883
rect 18325 11843 18383 11849
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 18785 11883 18843 11889
rect 18785 11849 18797 11883
rect 18831 11880 18843 11883
rect 18874 11880 18880 11892
rect 18831 11852 18880 11880
rect 18831 11849 18843 11852
rect 18785 11843 18843 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 20346 11880 20352 11892
rect 19996 11852 20352 11880
rect 8680 11812 8708 11840
rect 8326 11784 8708 11812
rect 8757 11815 8815 11821
rect 8757 11781 8769 11815
rect 8803 11812 8815 11815
rect 10321 11815 10379 11821
rect 8803 11784 9812 11812
rect 8803 11781 8815 11784
rect 8757 11775 8815 11781
rect 9508 11716 9674 11744
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11676 9091 11679
rect 9122 11676 9128 11688
rect 9079 11648 9128 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9508 11617 9536 11716
rect 9493 11611 9551 11617
rect 9493 11608 9505 11611
rect 8956 11580 9505 11608
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 8956 11540 8984 11580
rect 9493 11577 9505 11580
rect 9539 11577 9551 11611
rect 9646 11608 9674 11716
rect 9784 11676 9812 11784
rect 10321 11781 10333 11815
rect 10367 11812 10379 11815
rect 14366 11812 14372 11824
rect 10367 11784 14372 11812
rect 10367 11781 10379 11784
rect 10321 11775 10379 11781
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 14476 11784 15608 11812
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11744 11667 11747
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 11655 11716 12265 11744
rect 11655 11713 11667 11716
rect 11609 11707 11667 11713
rect 12253 11713 12265 11716
rect 12299 11744 12311 11747
rect 13449 11747 13507 11753
rect 12299 11716 12664 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 9784 11648 10425 11676
rect 10413 11645 10425 11648
rect 10459 11676 10471 11679
rect 11054 11676 11060 11688
rect 10459 11648 11060 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11940 11648 11989 11676
rect 11940 11636 11946 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 10226 11608 10232 11620
rect 9646 11580 10232 11608
rect 9493 11571 9551 11577
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 4028 11512 8984 11540
rect 9401 11543 9459 11549
rect 4028 11500 4034 11512
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9674 11540 9680 11552
rect 9447 11512 9680 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9674 11500 9680 11512
rect 9732 11540 9738 11552
rect 9858 11540 9864 11552
rect 9732 11512 9864 11540
rect 9732 11500 9738 11512
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 11333 11543 11391 11549
rect 11333 11509 11345 11543
rect 11379 11540 11391 11543
rect 11974 11540 11980 11552
rect 11379 11512 11980 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12636 11540 12664 11716
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 14476 11744 14504 11784
rect 13495 11716 14504 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 15580 11753 15608 11784
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 16666 11812 16672 11824
rect 16540 11784 16672 11812
rect 16540 11772 16546 11784
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 16758 11772 16764 11824
rect 16816 11812 16822 11824
rect 17586 11812 17592 11824
rect 16816 11784 17592 11812
rect 16816 11772 16822 11784
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 19794 11812 19800 11824
rect 18248 11784 19800 11812
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14608 11716 14657 11744
rect 14608 11704 14614 11716
rect 14645 11713 14657 11716
rect 14691 11744 14703 11747
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 14691 11716 15301 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 16776 11744 16804 11772
rect 15611 11716 16804 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 12802 11636 12808 11688
rect 12860 11676 12866 11688
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 12860 11648 13553 11676
rect 12860 11636 12866 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 13078 11568 13084 11620
rect 13136 11568 13142 11620
rect 13740 11608 13768 11639
rect 14734 11636 14740 11688
rect 14792 11636 14798 11688
rect 14826 11636 14832 11688
rect 14884 11636 14890 11688
rect 14844 11608 14872 11636
rect 13740 11580 14872 11608
rect 15304 11608 15332 11707
rect 17218 11704 17224 11756
rect 17276 11704 17282 11756
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 18248 11685 18276 11784
rect 19794 11772 19800 11784
rect 19852 11812 19858 11824
rect 19996 11812 20024 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 20772 11852 21189 11880
rect 20772 11840 20778 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 21450 11840 21456 11892
rect 21508 11840 21514 11892
rect 19852 11784 20024 11812
rect 19852 11772 19858 11784
rect 20070 11772 20076 11824
rect 20128 11812 20134 11824
rect 21545 11815 21603 11821
rect 21545 11812 21557 11815
rect 20128 11784 21557 11812
rect 20128 11772 20134 11784
rect 21545 11781 21557 11784
rect 21591 11812 21603 11815
rect 25958 11812 25964 11824
rect 21591 11784 25964 11812
rect 21591 11781 21603 11784
rect 21545 11775 21603 11781
rect 25958 11772 25964 11784
rect 26016 11772 26022 11824
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19426 11744 19432 11756
rect 19383 11716 19432 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20898 11744 20904 11756
rect 20404 11716 20904 11744
rect 20404 11704 20410 11716
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 24394 11744 24400 11756
rect 23523 11716 24400 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 25130 11704 25136 11756
rect 25188 11704 25194 11756
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 16540 11648 16957 11676
rect 16540 11636 16546 11648
rect 16945 11645 16957 11648
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20036 11648 20729 11676
rect 20036 11636 20042 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 23017 11679 23075 11685
rect 23017 11645 23029 11679
rect 23063 11645 23075 11679
rect 23017 11639 23075 11645
rect 17589 11611 17647 11617
rect 15304 11580 17540 11608
rect 14642 11540 14648 11552
rect 12636 11512 14648 11540
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16390 11540 16396 11552
rect 15344 11512 16396 11540
rect 15344 11500 15350 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 17512 11540 17540 11580
rect 17589 11577 17601 11611
rect 17635 11608 17647 11611
rect 21450 11608 21456 11620
rect 17635 11580 21456 11608
rect 17635 11577 17647 11580
rect 17589 11571 17647 11577
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 23032 11608 23060 11639
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 24854 11608 24860 11620
rect 23032 11580 24860 11608
rect 24854 11568 24860 11580
rect 24912 11568 24918 11620
rect 18598 11540 18604 11552
rect 17512 11512 18604 11540
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 19426 11500 19432 11552
rect 19484 11500 19490 11552
rect 20162 11500 20168 11552
rect 20220 11500 20226 11552
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 21818 11540 21824 11552
rect 20312 11512 21824 11540
rect 20312 11500 20318 11512
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 23290 11500 23296 11552
rect 23348 11540 23354 11552
rect 25774 11540 25780 11552
rect 23348 11512 25780 11540
rect 23348 11500 23354 11512
rect 25774 11500 25780 11512
rect 25832 11500 25838 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 12710 11296 12716 11348
rect 12768 11336 12774 11348
rect 12894 11336 12900 11348
rect 12768 11308 12900 11336
rect 12768 11296 12774 11308
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 15194 11336 15200 11348
rect 13044 11308 15200 11336
rect 13044 11296 13050 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 16356 11308 17233 11336
rect 16356 11296 16362 11308
rect 17221 11305 17233 11308
rect 17267 11336 17279 11339
rect 17267 11308 17816 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 10594 11228 10600 11280
rect 10652 11268 10658 11280
rect 10873 11271 10931 11277
rect 10873 11268 10885 11271
rect 10652 11240 10885 11268
rect 10652 11228 10658 11240
rect 10873 11237 10885 11240
rect 10919 11237 10931 11271
rect 10873 11231 10931 11237
rect 12161 11271 12219 11277
rect 12161 11237 12173 11271
rect 12207 11268 12219 11271
rect 12618 11268 12624 11280
rect 12207 11240 12624 11268
rect 12207 11237 12219 11240
rect 12161 11231 12219 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 13725 11271 13783 11277
rect 12912 11240 13676 11268
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 10410 11200 10416 11212
rect 9447 11172 10416 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 10410 11160 10416 11172
rect 10468 11200 10474 11212
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 10468 11172 11529 11200
rect 10468 11160 10474 11172
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11200 11759 11203
rect 12912 11200 12940 11240
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 11747 11172 12940 11200
rect 13004 11172 13185 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 13004 11132 13032 11172
rect 13173 11169 13185 11172
rect 13219 11200 13231 11203
rect 13538 11200 13544 11212
rect 13219 11172 13544 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 13648 11200 13676 11240
rect 13725 11237 13737 11271
rect 13771 11268 13783 11271
rect 13906 11268 13912 11280
rect 13771 11240 13912 11268
rect 13771 11237 13783 11240
rect 13725 11231 13783 11237
rect 13906 11228 13912 11240
rect 13964 11268 13970 11280
rect 14458 11268 14464 11280
rect 13964 11240 14464 11268
rect 13964 11228 13970 11240
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 16482 11228 16488 11280
rect 16540 11268 16546 11280
rect 16669 11271 16727 11277
rect 16669 11268 16681 11271
rect 16540 11240 16681 11268
rect 16540 11228 16546 11240
rect 16669 11237 16681 11240
rect 16715 11237 16727 11271
rect 16669 11231 16727 11237
rect 17034 11228 17040 11280
rect 17092 11268 17098 11280
rect 17310 11268 17316 11280
rect 17092 11240 17316 11268
rect 17092 11228 17098 11240
rect 17310 11228 17316 11240
rect 17368 11228 17374 11280
rect 17788 11268 17816 11308
rect 17862 11296 17868 11348
rect 17920 11296 17926 11348
rect 20254 11336 20260 11348
rect 18800 11308 20260 11336
rect 18800 11268 18828 11308
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20438 11336 20444 11348
rect 20395 11308 20444 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 20714 11296 20720 11348
rect 20772 11336 20778 11348
rect 22097 11339 22155 11345
rect 22097 11336 22109 11339
rect 20772 11308 22109 11336
rect 20772 11296 20778 11308
rect 22097 11305 22109 11308
rect 22143 11336 22155 11339
rect 23290 11336 23296 11348
rect 22143 11308 23296 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 24026 11296 24032 11348
rect 24084 11336 24090 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 24084 11308 25053 11336
rect 24084 11296 24090 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 17788 11240 18828 11268
rect 18877 11271 18935 11277
rect 18877 11237 18889 11271
rect 18923 11268 18935 11271
rect 20622 11268 20628 11280
rect 18923 11240 20628 11268
rect 18923 11237 18935 11240
rect 18877 11231 18935 11237
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 22738 11228 22744 11280
rect 22796 11268 22802 11280
rect 22796 11240 25268 11268
rect 22796 11228 22802 11240
rect 13817 11203 13875 11209
rect 13817 11200 13829 11203
rect 13648 11172 13829 11200
rect 13817 11169 13829 11172
rect 13863 11200 13875 11203
rect 14090 11200 14096 11212
rect 13863 11172 14096 11200
rect 13863 11169 13875 11172
rect 13817 11163 13875 11169
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 15930 11200 15936 11212
rect 14967 11172 15936 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 15930 11160 15936 11172
rect 15988 11200 15994 11212
rect 17402 11200 17408 11212
rect 15988 11172 17408 11200
rect 15988 11160 15994 11172
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 19334 11200 19340 11212
rect 18371 11172 19340 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19797 11203 19855 11209
rect 19797 11169 19809 11203
rect 19843 11200 19855 11203
rect 22646 11200 22652 11212
rect 19843 11172 22652 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 23290 11160 23296 11212
rect 23348 11160 23354 11212
rect 11112 11104 13032 11132
rect 13081 11135 13139 11141
rect 11112 11092 11118 11104
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 14826 11132 14832 11144
rect 13127 11104 14832 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 18782 11132 18788 11144
rect 18463 11104 18788 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 18782 11092 18788 11104
rect 18840 11132 18846 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18840 11104 19257 11132
rect 18840 11092 18846 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20772 11104 21005 11132
rect 20772 11092 20778 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 21508 11104 21557 11132
rect 21508 11092 21514 11104
rect 21545 11101 21557 11104
rect 21591 11101 21603 11135
rect 21545 11095 21603 11101
rect 24026 11092 24032 11144
rect 24084 11092 24090 11144
rect 25240 11141 25268 11240
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11101 25283 11135
rect 25225 11095 25283 11101
rect 10410 11024 10416 11076
rect 10468 11024 10474 11076
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 12584 11036 12664 11064
rect 12584 11024 12590 11036
rect 11790 10956 11796 11008
rect 11848 10956 11854 11008
rect 12636 11005 12664 11036
rect 12710 11024 12716 11076
rect 12768 11064 12774 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 12768 11036 14289 11064
rect 12768 11024 12774 11036
rect 14277 11033 14289 11036
rect 14323 11033 14335 11067
rect 14277 11027 14335 11033
rect 14458 11024 14464 11076
rect 14516 11064 14522 11076
rect 14516 11036 15056 11064
rect 14516 11024 14522 11036
rect 15028 11008 15056 11036
rect 15194 11024 15200 11076
rect 15252 11024 15258 11076
rect 16666 11064 16672 11076
rect 16422 11036 16672 11064
rect 16666 11024 16672 11036
rect 16724 11064 16730 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16724 11036 16957 11064
rect 16724 11024 16730 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 16945 11027 17003 11033
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17368 11036 17601 11064
rect 17368 11024 17374 11036
rect 17589 11033 17601 11036
rect 17635 11064 17647 11067
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 17635 11036 18521 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 18509 11027 18567 11033
rect 20806 11024 20812 11076
rect 20864 11024 20870 11076
rect 12621 10999 12679 11005
rect 12621 10965 12633 10999
rect 12667 10965 12679 10999
rect 12621 10959 12679 10965
rect 12986 10956 12992 11008
rect 13044 10956 13050 11008
rect 15010 10956 15016 11008
rect 15068 10956 15074 11008
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19852 10968 19901 10996
rect 19852 10956 19858 10968
rect 19889 10965 19901 10968
rect 19935 10965 19947 10999
rect 19889 10959 19947 10965
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 21450 10996 21456 11008
rect 20036 10968 21456 10996
rect 20036 10956 20042 10968
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 21726 10956 21732 11008
rect 21784 10956 21790 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 10042 10792 10048 10804
rect 9999 10764 10048 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 12618 10752 12624 10804
rect 12676 10752 12682 10804
rect 12710 10752 12716 10804
rect 12768 10752 12774 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 14182 10792 14188 10804
rect 13863 10764 14188 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 15470 10792 15476 10804
rect 14384 10764 15476 10792
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 7852 10696 8493 10724
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7852 10461 7880 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 9858 10724 9864 10736
rect 9706 10696 9864 10724
rect 8481 10687 8539 10693
rect 9858 10684 9864 10696
rect 9916 10724 9922 10736
rect 10410 10724 10416 10736
rect 9916 10696 10416 10724
rect 9916 10684 9922 10696
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 11882 10684 11888 10736
rect 11940 10724 11946 10736
rect 14384 10724 14412 10764
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 15562 10752 15568 10804
rect 15620 10752 15626 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16298 10792 16304 10804
rect 15979 10764 16304 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 17037 10795 17095 10801
rect 17037 10761 17049 10795
rect 17083 10792 17095 10795
rect 19978 10792 19984 10804
rect 17083 10764 19984 10792
rect 17083 10761 17095 10764
rect 17037 10755 17095 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20257 10795 20315 10801
rect 20257 10761 20269 10795
rect 20303 10792 20315 10795
rect 22186 10792 22192 10804
rect 20303 10764 22192 10792
rect 20303 10761 20315 10764
rect 20257 10755 20315 10761
rect 22186 10752 22192 10764
rect 22244 10752 22250 10804
rect 24118 10792 24124 10804
rect 22756 10764 24124 10792
rect 18322 10724 18328 10736
rect 11940 10696 14412 10724
rect 11940 10684 11946 10696
rect 14182 10616 14188 10668
rect 14240 10616 14246 10668
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7156 10424 7849 10452
rect 7156 10412 7162 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8220 10452 8248 10551
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 11241 10591 11299 10597
rect 11241 10588 11253 10591
rect 8536 10560 11253 10588
rect 8536 10548 8542 10560
rect 11241 10557 11253 10560
rect 11287 10588 11299 10591
rect 11790 10588 11796 10600
rect 11287 10560 11796 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 11882 10548 11888 10600
rect 11940 10548 11946 10600
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 12452 10520 12480 10551
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 13722 10588 13728 10600
rect 12952 10560 13728 10588
rect 12952 10548 12958 10560
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 13906 10548 13912 10600
rect 13964 10588 13970 10600
rect 14384 10597 14412 10696
rect 14476 10696 18328 10724
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 13964 10560 14289 10588
rect 13964 10548 13970 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 13449 10523 13507 10529
rect 13449 10520 13461 10523
rect 10652 10492 12480 10520
rect 12912 10492 13461 10520
rect 10652 10480 10658 10492
rect 9122 10452 9128 10464
rect 8220 10424 9128 10452
rect 7837 10415 7895 10421
rect 9122 10412 9128 10424
rect 9180 10452 9186 10464
rect 9582 10452 9588 10464
rect 9180 10424 9588 10452
rect 9180 10412 9186 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10962 10452 10968 10464
rect 10468 10424 10968 10452
rect 10468 10412 10474 10424
rect 10962 10412 10968 10424
rect 11020 10452 11026 10464
rect 12912 10452 12940 10492
rect 13449 10489 13461 10492
rect 13495 10489 13507 10523
rect 13449 10483 13507 10489
rect 11020 10424 12940 10452
rect 13081 10455 13139 10461
rect 11020 10412 11026 10424
rect 13081 10421 13093 10455
rect 13127 10452 13139 10455
rect 14476 10452 14504 10696
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 19610 10724 19616 10736
rect 18432 10696 19616 10724
rect 15470 10616 15476 10668
rect 15528 10656 15534 10668
rect 15528 10628 16160 10656
rect 15528 10616 15534 10628
rect 16132 10600 16160 10628
rect 16850 10616 16856 10668
rect 16908 10616 16914 10668
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 17828 10628 18245 10656
rect 17828 10616 17834 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 16022 10588 16028 10600
rect 15344 10560 16028 10588
rect 15344 10548 15350 10560
rect 16022 10548 16028 10560
rect 16080 10548 16086 10600
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 18432 10588 18460 10696
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 19978 10656 19984 10668
rect 19935 10628 19984 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 16224 10560 18460 10588
rect 13127 10424 14504 10452
rect 13127 10421 13139 10424
rect 13081 10415 13139 10421
rect 15286 10412 15292 10464
rect 15344 10412 15350 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 16224 10452 16252 10560
rect 17494 10480 17500 10532
rect 17552 10480 17558 10532
rect 18417 10523 18475 10529
rect 18417 10489 18429 10523
rect 18463 10520 18475 10523
rect 19076 10520 19104 10619
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22278 10656 22284 10668
rect 22235 10628 22284 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 19610 10548 19616 10600
rect 19668 10548 19674 10600
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 20438 10588 20444 10600
rect 19843 10560 20444 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 20680 10560 21189 10588
rect 20680 10548 20686 10560
rect 21177 10557 21189 10560
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21266 10548 21272 10600
rect 21324 10548 21330 10600
rect 21450 10548 21456 10600
rect 21508 10588 21514 10600
rect 22756 10588 22784 10764
rect 24118 10752 24124 10764
rect 24176 10752 24182 10804
rect 23382 10684 23388 10736
rect 23440 10684 23446 10736
rect 25133 10727 25191 10733
rect 25133 10724 25145 10727
rect 24610 10696 25145 10724
rect 25133 10693 25145 10696
rect 25179 10724 25191 10727
rect 25314 10724 25320 10736
rect 25179 10696 25320 10724
rect 25179 10693 25191 10696
rect 25133 10687 25191 10693
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 21508 10560 22784 10588
rect 21508 10548 21514 10560
rect 22830 10548 22836 10600
rect 22888 10588 22894 10600
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22888 10560 23121 10588
rect 22888 10548 22894 10560
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23109 10551 23167 10557
rect 20717 10523 20775 10529
rect 20717 10520 20729 10523
rect 18463 10492 19012 10520
rect 19076 10492 20729 10520
rect 18463 10489 18475 10492
rect 18417 10483 18475 10489
rect 15620 10424 16252 10452
rect 15620 10412 15626 10424
rect 18782 10412 18788 10464
rect 18840 10452 18846 10464
rect 18877 10455 18935 10461
rect 18877 10452 18889 10455
rect 18840 10424 18889 10452
rect 18840 10412 18846 10424
rect 18877 10421 18889 10424
rect 18923 10421 18935 10455
rect 18984 10452 19012 10492
rect 20717 10489 20729 10492
rect 20763 10489 20775 10523
rect 21284 10520 21312 10548
rect 21634 10520 21640 10532
rect 21284 10492 21640 10520
rect 20717 10483 20775 10489
rect 21634 10480 21640 10492
rect 21692 10480 21698 10532
rect 22094 10520 22100 10532
rect 21744 10492 22100 10520
rect 21744 10452 21772 10492
rect 22094 10480 22100 10492
rect 22152 10480 22158 10532
rect 18984 10424 21772 10452
rect 18877 10415 18935 10421
rect 22002 10412 22008 10464
rect 22060 10412 22066 10464
rect 22462 10412 22468 10464
rect 22520 10412 22526 10464
rect 22738 10412 22744 10464
rect 22796 10452 22802 10464
rect 23474 10452 23480 10464
rect 22796 10424 23480 10452
rect 22796 10412 22802 10424
rect 23474 10412 23480 10424
rect 23532 10412 23538 10464
rect 24118 10412 24124 10464
rect 24176 10452 24182 10464
rect 24857 10455 24915 10461
rect 24857 10452 24869 10455
rect 24176 10424 24869 10452
rect 24176 10412 24182 10424
rect 24857 10421 24869 10424
rect 24903 10421 24915 10455
rect 24857 10415 24915 10421
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 11606 10208 11612 10260
rect 11664 10208 11670 10260
rect 12406 10220 12940 10248
rect 12406 10180 12434 10220
rect 10612 10152 12434 10180
rect 12805 10183 12863 10189
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9582 10112 9588 10124
rect 9355 10084 9588 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10612 10112 10640 10152
rect 12805 10149 12817 10183
rect 12851 10149 12863 10183
rect 12912 10180 12940 10220
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 13780 10220 14565 10248
rect 13780 10208 13786 10220
rect 14553 10217 14565 10220
rect 14599 10217 14611 10251
rect 14553 10211 14611 10217
rect 15562 10208 15568 10260
rect 15620 10208 15626 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 19978 10248 19984 10260
rect 16080 10220 19984 10248
rect 16080 10208 16086 10220
rect 19978 10208 19984 10220
rect 20036 10248 20042 10260
rect 20165 10251 20223 10257
rect 20165 10248 20177 10251
rect 20036 10220 20177 10248
rect 20036 10208 20042 10220
rect 20165 10217 20177 10220
rect 20211 10217 20223 10251
rect 20165 10211 20223 10217
rect 24578 10208 24584 10260
rect 24636 10208 24642 10260
rect 12912 10152 13952 10180
rect 12805 10143 12863 10149
rect 10192 10084 10640 10112
rect 10192 10072 10198 10084
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12820 10112 12848 10143
rect 12400 10084 12848 10112
rect 13449 10115 13507 10121
rect 12400 10072 12406 10084
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13538 10112 13544 10124
rect 13495 10084 13544 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 11882 10004 11888 10056
rect 11940 10044 11946 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 11940 10016 13185 10044
rect 11940 10004 11946 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 9306 9936 9312 9988
rect 9364 9976 9370 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9364 9948 9597 9976
rect 9364 9936 9370 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 10962 9976 10968 9988
rect 10810 9948 10968 9976
rect 9585 9939 9643 9945
rect 10962 9936 10968 9948
rect 11020 9976 11026 9988
rect 11606 9976 11612 9988
rect 11020 9948 11612 9976
rect 11020 9936 11026 9948
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 11977 9979 12035 9985
rect 11977 9945 11989 9979
rect 12023 9976 12035 9979
rect 13722 9976 13728 9988
rect 12023 9948 13728 9976
rect 12023 9945 12035 9948
rect 11977 9939 12035 9945
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 13924 9985 13952 10152
rect 14182 10140 14188 10192
rect 14240 10180 14246 10192
rect 16574 10180 16580 10192
rect 14240 10152 16580 10180
rect 14240 10140 14246 10152
rect 16574 10140 16580 10152
rect 16632 10180 16638 10192
rect 20530 10180 20536 10192
rect 16632 10152 20536 10180
rect 16632 10140 16638 10152
rect 20530 10140 20536 10152
rect 20588 10140 20594 10192
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 14458 10112 14464 10124
rect 14323 10084 14464 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 14458 10072 14464 10084
rect 14516 10112 14522 10124
rect 15102 10112 15108 10124
rect 14516 10084 15108 10112
rect 14516 10072 14522 10084
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 16776 10084 18368 10112
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 16776 10044 16804 10084
rect 14792 10016 16804 10044
rect 16853 10047 16911 10053
rect 14792 10004 14798 10016
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 17678 10044 17684 10056
rect 16899 10016 17684 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 13909 9979 13967 9985
rect 13909 9945 13921 9979
rect 13955 9976 13967 9979
rect 15013 9979 15071 9985
rect 15013 9976 15025 9979
rect 13955 9948 15025 9976
rect 13955 9945 13967 9948
rect 13909 9939 13967 9945
rect 15013 9945 15025 9948
rect 15059 9976 15071 9979
rect 17862 9976 17868 9988
rect 15059 9948 17868 9976
rect 15059 9945 15071 9948
rect 15013 9939 15071 9945
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 18340 9985 18368 10084
rect 18414 10072 18420 10124
rect 18472 10072 18478 10124
rect 18598 10072 18604 10124
rect 18656 10072 18662 10124
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 20809 10115 20867 10121
rect 20809 10112 20821 10115
rect 19392 10084 20821 10112
rect 19392 10072 19398 10084
rect 20809 10081 20821 10084
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 20898 10072 20904 10124
rect 20956 10112 20962 10124
rect 21358 10112 21364 10124
rect 20956 10084 21364 10112
rect 20956 10072 20962 10084
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 21542 10072 21548 10124
rect 21600 10112 21606 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 21600 10084 23305 10112
rect 21600 10072 21606 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23385 10115 23443 10121
rect 23385 10081 23397 10115
rect 23431 10112 23443 10115
rect 24118 10112 24124 10124
rect 23431 10084 24124 10112
rect 23431 10081 23443 10084
rect 23385 10075 23443 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 18325 9979 18383 9985
rect 18325 9945 18337 9979
rect 18371 9945 18383 9979
rect 18432 9976 18460 10072
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 19024 10016 20545 10044
rect 19024 10004 19030 10016
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 22612 10016 24777 10044
rect 22612 10004 22618 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 19061 9979 19119 9985
rect 19061 9976 19073 9979
rect 18432 9948 19073 9976
rect 18325 9939 18383 9945
rect 19061 9945 19073 9948
rect 19107 9945 19119 9979
rect 19061 9939 19119 9945
rect 19613 9979 19671 9985
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 20254 9976 20260 9988
rect 19659 9948 20260 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 20254 9936 20260 9948
rect 20312 9936 20318 9988
rect 21358 9936 21364 9988
rect 21416 9936 21422 9988
rect 22186 9936 22192 9988
rect 22244 9976 22250 9988
rect 25038 9976 25044 9988
rect 22244 9948 25044 9976
rect 22244 9936 22250 9948
rect 25038 9936 25044 9948
rect 25096 9936 25102 9988
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 12802 9908 12808 9920
rect 12115 9880 12808 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 13446 9908 13452 9920
rect 13311 9880 13452 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9908 14979 9911
rect 15470 9908 15476 9920
rect 14967 9880 15476 9908
rect 14967 9877 14979 9880
rect 14921 9871 14979 9877
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 15841 9911 15899 9917
rect 15841 9908 15853 9911
rect 15620 9880 15853 9908
rect 15620 9868 15626 9880
rect 15841 9877 15853 9880
rect 15887 9908 15899 9911
rect 16022 9908 16028 9920
rect 15887 9880 16028 9908
rect 15887 9877 15899 9880
rect 15841 9871 15899 9877
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 16301 9911 16359 9917
rect 16301 9877 16313 9911
rect 16347 9908 16359 9911
rect 16390 9908 16396 9920
rect 16347 9880 16396 9908
rect 16347 9877 16359 9880
rect 16301 9871 16359 9877
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16816 9880 16957 9908
rect 16816 9868 16822 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 17957 9911 18015 9917
rect 17957 9877 17969 9911
rect 18003 9908 18015 9911
rect 18230 9908 18236 9920
rect 18003 9880 18236 9908
rect 18003 9877 18015 9880
rect 17957 9871 18015 9877
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 19518 9868 19524 9920
rect 19576 9868 19582 9920
rect 19794 9868 19800 9920
rect 19852 9908 19858 9920
rect 19978 9908 19984 9920
rect 19852 9880 19984 9908
rect 19852 9868 19858 9880
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 21634 9868 21640 9920
rect 21692 9908 21698 9920
rect 22281 9911 22339 9917
rect 22281 9908 22293 9911
rect 21692 9880 22293 9908
rect 21692 9868 21698 9880
rect 22281 9877 22293 9880
rect 22327 9877 22339 9911
rect 22281 9871 22339 9877
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 22833 9911 22891 9917
rect 22833 9908 22845 9911
rect 22428 9880 22845 9908
rect 22428 9868 22434 9880
rect 22833 9877 22845 9880
rect 22879 9877 22891 9911
rect 22833 9871 22891 9877
rect 23201 9911 23259 9917
rect 23201 9877 23213 9911
rect 23247 9908 23259 9911
rect 24578 9908 24584 9920
rect 23247 9880 24584 9908
rect 23247 9877 23259 9880
rect 23201 9871 23259 9877
rect 24578 9868 24584 9880
rect 24636 9868 24642 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 12342 9704 12348 9716
rect 7156 9676 12348 9704
rect 7156 9664 7162 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15470 9704 15476 9716
rect 15344 9676 15476 9704
rect 15344 9664 15350 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 18966 9704 18972 9716
rect 17460 9676 18972 9704
rect 17460 9664 17466 9676
rect 18966 9664 18972 9676
rect 19024 9704 19030 9716
rect 20898 9704 20904 9716
rect 19024 9676 19104 9704
rect 19024 9664 19030 9676
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 8846 9636 8852 9648
rect 3936 9608 8852 9636
rect 3936 9596 3942 9608
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 11664 9608 12466 9636
rect 11664 9596 11670 9608
rect 16114 9596 16120 9648
rect 16172 9636 16178 9648
rect 16298 9636 16304 9648
rect 16172 9608 16304 9636
rect 16172 9596 16178 9608
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 16942 9636 16948 9648
rect 16724 9608 16948 9636
rect 16724 9596 16730 9608
rect 16942 9596 16948 9608
rect 17000 9636 17006 9648
rect 17000 9622 17618 9636
rect 17000 9608 17632 9622
rect 17000 9596 17006 9608
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 15378 9568 15384 9580
rect 14323 9540 15384 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9537 15531 9571
rect 17310 9568 17316 9580
rect 15473 9531 15531 9537
rect 15672 9540 17316 9568
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 11514 9500 11520 9512
rect 10744 9472 11520 9500
rect 10744 9460 10750 9472
rect 11514 9460 11520 9472
rect 11572 9500 11578 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11572 9472 11713 9500
rect 11572 9460 11578 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12710 9500 12716 9512
rect 12023 9472 12716 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 13814 9500 13820 9512
rect 13495 9472 13820 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14366 9500 14372 9512
rect 14056 9472 14372 9500
rect 14056 9460 14062 9472
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 13780 9404 13921 9432
rect 13780 9392 13786 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 14826 9392 14832 9444
rect 14884 9432 14890 9444
rect 15105 9435 15163 9441
rect 15105 9432 15117 9435
rect 14884 9404 15117 9432
rect 14884 9392 14890 9404
rect 15105 9401 15117 9404
rect 15151 9401 15163 9435
rect 15488 9432 15516 9531
rect 15672 9512 15700 9540
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15654 9500 15660 9512
rect 15611 9472 15660 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 15838 9500 15844 9512
rect 15795 9472 15844 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16080 9472 16957 9500
rect 16080 9460 16086 9472
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 17604 9500 17632 9608
rect 18690 9596 18696 9648
rect 18748 9636 18754 9648
rect 18785 9639 18843 9645
rect 18785 9636 18797 9639
rect 18748 9608 18797 9636
rect 18748 9596 18754 9608
rect 18785 9605 18797 9608
rect 18831 9605 18843 9639
rect 18785 9599 18843 9605
rect 19076 9577 19104 9676
rect 20640 9676 20904 9704
rect 19794 9596 19800 9648
rect 19852 9636 19858 9648
rect 20640 9636 20668 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 22005 9707 22063 9713
rect 22005 9704 22017 9707
rect 21140 9676 22017 9704
rect 21140 9664 21146 9676
rect 22005 9673 22017 9676
rect 22051 9673 22063 9707
rect 23382 9704 23388 9716
rect 22005 9667 22063 9673
rect 22848 9676 23388 9704
rect 19852 9608 20668 9636
rect 19852 9596 19858 9608
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 21450 9636 21456 9648
rect 20772 9608 21456 9636
rect 20772 9596 20778 9608
rect 21450 9596 21456 9608
rect 21508 9596 21514 9648
rect 21542 9596 21548 9648
rect 21600 9636 21606 9648
rect 22738 9636 22744 9648
rect 21600 9608 22744 9636
rect 21600 9596 21606 9608
rect 22738 9596 22744 9608
rect 22796 9636 22802 9648
rect 22848 9636 22876 9676
rect 23382 9664 23388 9676
rect 23440 9704 23446 9716
rect 25314 9704 25320 9716
rect 23440 9676 25320 9704
rect 23440 9664 23446 9676
rect 25314 9664 25320 9676
rect 25372 9664 25378 9716
rect 22796 9608 22876 9636
rect 22796 9596 22802 9608
rect 23474 9596 23480 9648
rect 23532 9596 23538 9648
rect 24118 9596 24124 9648
rect 24176 9596 24182 9648
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 19300 9540 20085 9568
rect 19300 9528 19306 9540
rect 20073 9537 20085 9540
rect 20119 9537 20131 9571
rect 20073 9531 20131 9537
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 22554 9568 22560 9580
rect 21315 9540 22560 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 22554 9528 22560 9540
rect 22612 9528 22618 9580
rect 24946 9528 24952 9580
rect 25004 9568 25010 9580
rect 25041 9571 25099 9577
rect 25041 9568 25053 9571
rect 25004 9540 25053 9568
rect 25004 9528 25010 9540
rect 25041 9537 25053 9540
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 17604 9472 19334 9500
rect 16945 9463 17003 9469
rect 15488 9404 16436 9432
rect 15105 9395 15163 9401
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9364 11391 9367
rect 11514 9364 11520 9376
rect 11379 9336 11520 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 16408 9373 16436 9404
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 17034 9432 17040 9444
rect 16632 9404 17040 9432
rect 16632 9392 16638 9404
rect 17034 9392 17040 9404
rect 17092 9432 17098 9444
rect 17313 9435 17371 9441
rect 17313 9432 17325 9435
rect 17092 9404 17325 9432
rect 17092 9392 17098 9404
rect 17313 9401 17325 9404
rect 17359 9401 17371 9435
rect 19306 9432 19334 9472
rect 22646 9460 22652 9512
rect 22704 9460 22710 9512
rect 24397 9503 24455 9509
rect 24397 9469 24409 9503
rect 24443 9469 24455 9503
rect 24397 9463 24455 9469
rect 19429 9435 19487 9441
rect 19429 9432 19441 9435
rect 19306 9404 19441 9432
rect 17313 9395 17371 9401
rect 19429 9401 19441 9404
rect 19475 9432 19487 9435
rect 19794 9432 19800 9444
rect 19475 9404 19800 9432
rect 19475 9401 19487 9404
rect 19429 9395 19487 9401
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 22830 9432 22836 9444
rect 22152 9404 22836 9432
rect 22152 9392 22158 9404
rect 22830 9392 22836 9404
rect 22888 9432 22894 9444
rect 22888 9404 23152 9432
rect 22888 9392 22894 9404
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 14424 9336 16129 9364
rect 14424 9324 14430 9336
rect 16117 9333 16129 9336
rect 16163 9333 16175 9367
rect 16117 9327 16175 9333
rect 16393 9367 16451 9373
rect 16393 9333 16405 9367
rect 16439 9364 16451 9367
rect 16666 9364 16672 9376
rect 16439 9336 16672 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16853 9367 16911 9373
rect 16853 9333 16865 9367
rect 16899 9364 16911 9367
rect 17402 9364 17408 9376
rect 16899 9336 17408 9364
rect 16899 9333 16911 9336
rect 16853 9327 16911 9333
rect 17402 9324 17408 9336
rect 17460 9364 17466 9376
rect 21358 9364 21364 9376
rect 17460 9336 21364 9364
rect 17460 9324 17466 9336
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 23124 9364 23152 9404
rect 24412 9364 24440 9463
rect 23124 9336 24440 9364
rect 24854 9324 24860 9376
rect 24912 9324 24918 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12618 9160 12624 9172
rect 12400 9132 12624 9160
rect 12400 9120 12406 9132
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 12860 9132 14289 9160
rect 12860 9120 12866 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 15933 9163 15991 9169
rect 15933 9160 15945 9163
rect 15804 9132 15945 9160
rect 15804 9120 15810 9132
rect 15933 9129 15945 9132
rect 15979 9129 15991 9163
rect 15933 9123 15991 9129
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 17954 9160 17960 9172
rect 16724 9132 17960 9160
rect 16724 9120 16730 9132
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 19613 9163 19671 9169
rect 19613 9160 19625 9163
rect 19392 9132 19625 9160
rect 19392 9120 19398 9132
rect 19613 9129 19625 9132
rect 19659 9129 19671 9163
rect 19613 9123 19671 9129
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 12492 9064 13001 9092
rect 12492 9052 12498 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 12989 9055 13047 9061
rect 13998 9052 14004 9104
rect 14056 9092 14062 9104
rect 15473 9095 15531 9101
rect 15473 9092 15485 9095
rect 14056 9064 15485 9092
rect 14056 9052 14062 9064
rect 15473 9061 15485 9064
rect 15519 9092 15531 9095
rect 15654 9092 15660 9104
rect 15519 9064 15660 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17129 9095 17187 9101
rect 17129 9092 17141 9095
rect 17092 9064 17141 9092
rect 17092 9052 17098 9064
rect 17129 9061 17141 9064
rect 17175 9061 17187 9095
rect 19978 9092 19984 9104
rect 17129 9055 17187 9061
rect 17880 9064 19984 9092
rect 10594 8984 10600 9036
rect 10652 8984 10658 9036
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 14516 8996 14841 9024
rect 14516 8984 14522 8996
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16356 8996 16497 9024
rect 16356 8984 16362 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 17678 8984 17684 9036
rect 17736 8984 17742 9036
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 10166 8860 10548 8888
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9306 8820 9312 8832
rect 9171 8792 9312 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 10520 8820 10548 8860
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10888 8888 10916 8919
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 12676 8928 12725 8956
rect 12676 8916 12682 8928
rect 12713 8925 12725 8928
rect 12759 8956 12771 8959
rect 14476 8956 14504 8984
rect 12759 8928 14504 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 16022 8916 16028 8968
rect 16080 8956 16086 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 16080 8952 16252 8956
rect 16316 8952 17601 8956
rect 16080 8928 17601 8952
rect 16080 8916 16086 8928
rect 16224 8924 16344 8928
rect 17589 8925 17601 8928
rect 17635 8956 17647 8959
rect 17880 8956 17908 9064
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 19058 9024 19064 9036
rect 18012 8996 19064 9024
rect 18012 8984 18018 8996
rect 19058 8984 19064 8996
rect 19116 9024 19122 9036
rect 20990 9024 20996 9036
rect 19116 8996 20996 9024
rect 19116 8984 19122 8996
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 21361 9027 21419 9033
rect 21361 8993 21373 9027
rect 21407 9024 21419 9027
rect 22094 9024 22100 9036
rect 21407 8996 22100 9024
rect 21407 8993 21419 8996
rect 21361 8987 21419 8993
rect 22094 8984 22100 8996
rect 22152 8984 22158 9036
rect 25041 9027 25099 9033
rect 25041 9024 25053 9027
rect 22848 8996 25053 9024
rect 17635 8928 17908 8956
rect 18693 8959 18751 8965
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 19150 8956 19156 8968
rect 18739 8928 19156 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 22848 8965 22876 8996
rect 25041 8993 25053 8996
rect 25087 8993 25099 9027
rect 25041 8987 25099 8993
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21508 8928 22017 8956
rect 21508 8916 21514 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 10744 8860 10916 8888
rect 13357 8891 13415 8897
rect 10744 8848 10750 8860
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 13538 8888 13544 8900
rect 13403 8860 13544 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 13872 8860 14749 8888
rect 13872 8848 13878 8860
rect 14737 8857 14749 8860
rect 14783 8888 14795 8891
rect 14826 8888 14832 8900
rect 14783 8860 14832 8888
rect 14783 8857 14795 8860
rect 14737 8851 14795 8857
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 16393 8891 16451 8897
rect 16393 8888 16405 8891
rect 16224 8860 16405 8888
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 10520 8792 11253 8820
rect 11241 8789 11253 8792
rect 11287 8820 11299 8823
rect 11514 8820 11520 8832
rect 11287 8792 11520 8820
rect 11287 8789 11299 8792
rect 11241 8783 11299 8789
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 13449 8823 13507 8829
rect 13449 8789 13461 8823
rect 13495 8820 13507 8823
rect 14182 8820 14188 8832
rect 13495 8792 14188 8820
rect 13495 8789 13507 8792
rect 13449 8783 13507 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 14608 8792 14657 8820
rect 14608 8780 14614 8792
rect 14645 8789 14657 8792
rect 14691 8820 14703 8823
rect 15286 8820 15292 8832
rect 14691 8792 15292 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15378 8780 15384 8832
rect 15436 8780 15442 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16224 8820 16252 8860
rect 16393 8857 16405 8860
rect 16439 8857 16451 8891
rect 16393 8851 16451 8857
rect 17497 8891 17555 8897
rect 17497 8857 17509 8891
rect 17543 8857 17555 8891
rect 17497 8851 17555 8857
rect 15620 8792 16252 8820
rect 16301 8823 16359 8829
rect 15620 8780 15626 8792
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 17402 8820 17408 8832
rect 16347 8792 17408 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 17402 8780 17408 8792
rect 17460 8780 17466 8832
rect 17512 8820 17540 8851
rect 17862 8848 17868 8900
rect 17920 8888 17926 8900
rect 18414 8888 18420 8900
rect 17920 8860 18420 8888
rect 17920 8848 17926 8860
rect 18414 8848 18420 8860
rect 18472 8848 18478 8900
rect 18877 8891 18935 8897
rect 18877 8857 18889 8891
rect 18923 8888 18935 8891
rect 19518 8888 19524 8900
rect 18923 8860 19524 8888
rect 18923 8857 18935 8860
rect 18877 8851 18935 8857
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 19794 8848 19800 8900
rect 19852 8888 19858 8900
rect 21085 8891 21143 8897
rect 19852 8860 19918 8888
rect 19852 8848 19858 8860
rect 21085 8857 21097 8891
rect 21131 8857 21143 8891
rect 21085 8851 21143 8857
rect 18233 8823 18291 8829
rect 18233 8820 18245 8823
rect 17512 8792 18245 8820
rect 18233 8789 18245 8792
rect 18279 8820 18291 8823
rect 20346 8820 20352 8832
rect 18279 8792 20352 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 21100 8820 21128 8851
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 22848 8888 22876 8919
rect 24210 8916 24216 8968
rect 24268 8956 24274 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24268 8928 24593 8956
rect 24268 8916 24274 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 21232 8860 22876 8888
rect 23845 8891 23903 8897
rect 21232 8848 21238 8860
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 21266 8820 21272 8832
rect 21100 8792 21272 8820
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 21821 8823 21879 8829
rect 21821 8789 21833 8823
rect 21867 8820 21879 8823
rect 22186 8820 22192 8832
rect 21867 8792 22192 8820
rect 21867 8789 21879 8792
rect 21821 8783 21879 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 22373 8823 22431 8829
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 23382 8820 23388 8832
rect 22419 8792 23388 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 24762 8780 24768 8832
rect 24820 8780 24826 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 13354 8616 13360 8628
rect 12943 8588 13360 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 13354 8576 13360 8588
rect 13412 8616 13418 8628
rect 13412 8588 13952 8616
rect 13412 8576 13418 8588
rect 13924 8557 13952 8588
rect 14090 8576 14096 8628
rect 14148 8616 14154 8628
rect 21174 8616 21180 8628
rect 14148 8588 21180 8616
rect 14148 8576 14154 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 14458 8508 14464 8560
rect 14516 8508 14522 8560
rect 15396 8520 23980 8548
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 15010 8480 15016 8492
rect 14424 8452 15016 8480
rect 14424 8440 14430 8452
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 15396 8489 15424 8520
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 15381 8443 15439 8449
rect 15488 8452 17233 8480
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 13354 8372 13360 8424
rect 13412 8372 13418 8424
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 15488 8412 15516 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17862 8480 17868 8492
rect 17368 8452 17868 8480
rect 17368 8440 17374 8452
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18414 8440 18420 8492
rect 18472 8440 18478 8492
rect 18524 8452 20760 8480
rect 13964 8384 15516 8412
rect 13964 8372 13970 8384
rect 15654 8372 15660 8424
rect 15712 8372 15718 8424
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 17034 8372 17040 8424
rect 17092 8372 17098 8424
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 17328 8412 17356 8440
rect 18524 8412 18552 8452
rect 17175 8384 17356 8412
rect 17420 8384 18552 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8344 14151 8347
rect 14826 8344 14832 8356
rect 14139 8316 14832 8344
rect 14139 8313 14151 8316
rect 14093 8307 14151 8313
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 17420 8344 17448 8384
rect 19058 8372 19064 8424
rect 19116 8372 19122 8424
rect 20438 8372 20444 8424
rect 20496 8372 20502 8424
rect 15436 8316 17448 8344
rect 17589 8347 17647 8353
rect 15436 8304 15442 8316
rect 17589 8313 17601 8347
rect 17635 8344 17647 8347
rect 20622 8344 20628 8356
rect 17635 8316 20628 8344
rect 17635 8313 17647 8316
rect 17589 8307 17647 8313
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 20732 8344 20760 8452
rect 21450 8440 21456 8492
rect 21508 8440 21514 8492
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 23952 8489 23980 8520
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 22281 8483 22339 8489
rect 22281 8480 22293 8483
rect 22244 8452 22293 8480
rect 22244 8440 22250 8452
rect 22281 8449 22293 8452
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 22462 8372 22468 8424
rect 22520 8412 22526 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 22520 8384 22569 8412
rect 22520 8372 22526 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 21542 8344 21548 8356
rect 20732 8316 21548 8344
rect 21542 8304 21548 8316
rect 21600 8304 21606 8356
rect 21818 8304 21824 8356
rect 21876 8344 21882 8356
rect 24118 8344 24124 8356
rect 21876 8316 24124 8344
rect 21876 8304 21882 8316
rect 24118 8304 24124 8316
rect 24176 8304 24182 8356
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 22002 8276 22008 8288
rect 16264 8248 22008 8276
rect 16264 8236 16270 8248
rect 22002 8236 22008 8248
rect 22060 8276 22066 8288
rect 24486 8276 24492 8288
rect 22060 8248 24492 8276
rect 22060 8236 22066 8248
rect 24486 8236 24492 8248
rect 24544 8236 24550 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 14090 8072 14096 8084
rect 10376 8044 14096 8072
rect 10376 8032 10382 8044
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 15841 8075 15899 8081
rect 15841 8072 15853 8075
rect 14240 8044 15853 8072
rect 14240 8032 14246 8044
rect 15841 8041 15853 8044
rect 15887 8041 15899 8075
rect 25314 8072 25320 8084
rect 15841 8035 15899 8041
rect 18432 8044 25320 8072
rect 11790 7964 11796 8016
rect 11848 7964 11854 8016
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 15013 8007 15071 8013
rect 12768 7976 14412 8004
rect 12768 7964 12774 7976
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11882 7936 11888 7948
rect 11287 7908 11888 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 14384 7945 14412 7976
rect 15013 7973 15025 8007
rect 15059 8004 15071 8007
rect 17770 8004 17776 8016
rect 15059 7976 17776 8004
rect 15059 7973 15071 7976
rect 15013 7967 15071 7973
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 14369 7939 14427 7945
rect 13219 7908 14320 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11698 7868 11704 7880
rect 11471 7840 11704 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 14292 7868 14320 7908
rect 14369 7905 14381 7939
rect 14415 7905 14427 7939
rect 15194 7936 15200 7948
rect 14369 7899 14427 7905
rect 14568 7908 15200 7936
rect 14568 7868 14596 7908
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 15896 7908 16405 7936
rect 15896 7896 15902 7908
rect 16393 7905 16405 7908
rect 16439 7936 16451 7939
rect 17678 7936 17684 7948
rect 16439 7908 17684 7936
rect 16439 7905 16451 7908
rect 16393 7899 16451 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 18432 7945 18460 8044
rect 25314 8032 25320 8044
rect 25372 8032 25378 8084
rect 23474 7964 23480 8016
rect 23532 8004 23538 8016
rect 23845 8007 23903 8013
rect 23845 8004 23857 8007
rect 23532 7976 23857 8004
rect 23532 7964 23538 7976
rect 23845 7973 23857 7976
rect 23891 7973 23903 8007
rect 23845 7967 23903 7973
rect 24026 7964 24032 8016
rect 24084 8004 24090 8016
rect 24581 8007 24639 8013
rect 24581 8004 24593 8007
rect 24084 7976 24593 8004
rect 24084 7964 24090 7976
rect 24581 7973 24593 7976
rect 24627 7973 24639 8007
rect 24581 7967 24639 7973
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7905 18475 7939
rect 18417 7899 18475 7905
rect 21177 7939 21235 7945
rect 21177 7905 21189 7939
rect 21223 7905 21235 7939
rect 21177 7899 21235 7905
rect 22373 7939 22431 7945
rect 22373 7905 22385 7939
rect 22419 7936 22431 7939
rect 22830 7936 22836 7948
rect 22419 7908 22836 7936
rect 22419 7905 22431 7908
rect 22373 7899 22431 7905
rect 14292 7840 14596 7868
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 16114 7868 16120 7880
rect 14691 7840 16120 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 17218 7868 17224 7880
rect 16224 7840 17224 7868
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 8628 7772 13277 7800
rect 8628 7760 8634 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 16224 7800 16252 7840
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 20070 7868 20076 7880
rect 18923 7840 20076 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 13265 7763 13323 7769
rect 13740 7772 16252 7800
rect 11330 7692 11336 7744
rect 11388 7692 11394 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 12618 7732 12624 7744
rect 12575 7704 12624 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13740 7741 13768 7772
rect 16298 7760 16304 7812
rect 16356 7760 16362 7812
rect 16390 7760 16396 7812
rect 16448 7800 16454 7812
rect 21082 7800 21088 7812
rect 16448 7772 21088 7800
rect 16448 7760 16454 7772
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7701 13783 7735
rect 13725 7695 13783 7701
rect 14550 7692 14556 7744
rect 14608 7692 14614 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15381 7735 15439 7741
rect 15381 7732 15393 7735
rect 15344 7704 15393 7732
rect 15344 7692 15350 7704
rect 15381 7701 15393 7704
rect 15427 7732 15439 7735
rect 15838 7732 15844 7744
rect 15427 7704 15844 7732
rect 15427 7701 15439 7704
rect 15381 7695 15439 7701
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 16206 7692 16212 7744
rect 16264 7692 16270 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 19392 7704 19441 7732
rect 19392 7692 19398 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 19794 7692 19800 7744
rect 19852 7732 19858 7744
rect 19889 7735 19947 7741
rect 19889 7732 19901 7735
rect 19852 7704 19901 7732
rect 19852 7692 19858 7704
rect 19889 7701 19901 7704
rect 19935 7701 19947 7735
rect 21192 7732 21220 7899
rect 22830 7896 22836 7908
rect 22888 7896 22894 7948
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7868 21695 7871
rect 21818 7868 21824 7880
rect 21683 7840 21824 7868
rect 21683 7837 21695 7840
rect 21637 7831 21695 7837
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22094 7828 22100 7880
rect 22152 7828 22158 7880
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 23440 7854 23506 7868
rect 23440 7840 23520 7854
rect 23440 7828 23446 7840
rect 22554 7732 22560 7744
rect 21192 7704 22560 7732
rect 19889 7695 19947 7701
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 23492 7732 23520 7840
rect 23658 7760 23664 7812
rect 23716 7800 23722 7812
rect 24765 7803 24823 7809
rect 24765 7800 24777 7803
rect 23716 7772 24777 7800
rect 23716 7760 23722 7772
rect 24765 7769 24777 7772
rect 24811 7769 24823 7803
rect 24765 7763 24823 7769
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 23492 7704 24225 7732
rect 24213 7701 24225 7704
rect 24259 7732 24271 7735
rect 24670 7732 24676 7744
rect 24259 7704 24676 7732
rect 24259 7701 24271 7704
rect 24213 7695 24271 7701
rect 24670 7692 24676 7704
rect 24728 7692 24734 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 16850 7528 16856 7540
rect 13035 7500 16856 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17773 7531 17831 7537
rect 17773 7497 17785 7531
rect 17819 7528 17831 7531
rect 18322 7528 18328 7540
rect 17819 7500 18328 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 18690 7528 18696 7540
rect 18555 7500 18696 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 9582 7460 9588 7472
rect 9048 7432 9588 7460
rect 9048 7401 9076 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 11514 7460 11520 7472
rect 10534 7432 11520 7460
rect 11514 7420 11520 7432
rect 11572 7420 11578 7472
rect 14458 7420 14464 7472
rect 14516 7420 14522 7472
rect 15197 7463 15255 7469
rect 15197 7429 15209 7463
rect 15243 7460 15255 7463
rect 16482 7460 16488 7472
rect 15243 7432 16488 7460
rect 15243 7429 15255 7432
rect 15197 7423 15255 7429
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 16761 7463 16819 7469
rect 16761 7429 16773 7463
rect 16807 7460 16819 7463
rect 16942 7460 16948 7472
rect 16807 7432 16948 7460
rect 16807 7429 16819 7432
rect 16761 7423 16819 7429
rect 16942 7420 16948 7432
rect 17000 7460 17006 7472
rect 17862 7460 17868 7472
rect 17000 7432 17868 7460
rect 17000 7420 17006 7432
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 13814 7392 13820 7404
rect 12124 7364 13820 7392
rect 12124 7352 12130 7364
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 17681 7395 17739 7401
rect 16163 7364 16197 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 17727 7364 17908 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 10796 7296 12357 7324
rect 10796 7200 10824 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12526 7284 12532 7336
rect 12584 7284 12590 7336
rect 15102 7284 15108 7336
rect 15160 7324 15166 7336
rect 15473 7327 15531 7333
rect 15160 7296 15424 7324
rect 15160 7284 15166 7296
rect 11149 7259 11207 7265
rect 11149 7225 11161 7259
rect 11195 7256 11207 7259
rect 11514 7256 11520 7268
rect 11195 7228 11520 7256
rect 11195 7225 11207 7228
rect 11149 7219 11207 7225
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 11882 7216 11888 7268
rect 11940 7256 11946 7268
rect 15396 7256 15424 7296
rect 15473 7293 15485 7327
rect 15519 7324 15531 7327
rect 15930 7324 15936 7336
rect 15519 7296 15936 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16132 7324 16160 7355
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 16040 7296 16865 7324
rect 16040 7256 16068 7296
rect 16853 7293 16865 7296
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 11940 7228 14228 7256
rect 15396 7228 16068 7256
rect 16301 7259 16359 7265
rect 11940 7216 11946 7228
rect 10778 7148 10784 7200
rect 10836 7148 10842 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11422 7188 11428 7200
rect 11379 7160 11428 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 13596 7160 13737 7188
rect 13596 7148 13602 7160
rect 13725 7157 13737 7160
rect 13771 7157 13783 7191
rect 14200 7188 14228 7228
rect 16301 7225 16313 7259
rect 16347 7256 16359 7259
rect 17402 7256 17408 7268
rect 16347 7228 17408 7256
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 17402 7216 17408 7228
rect 17460 7216 17466 7268
rect 16574 7188 16580 7200
rect 14200 7160 16580 7188
rect 13725 7151 13783 7157
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16942 7148 16948 7200
rect 17000 7188 17006 7200
rect 17313 7191 17371 7197
rect 17313 7188 17325 7191
rect 17000 7160 17325 7188
rect 17000 7148 17006 7160
rect 17313 7157 17325 7160
rect 17359 7157 17371 7191
rect 17880 7188 17908 7364
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7324 18015 7327
rect 18524 7324 18552 7491
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19794 7488 19800 7540
rect 19852 7488 19858 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 20680 7500 21189 7528
rect 20680 7488 20686 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 19812 7460 19840 7488
rect 20530 7460 20536 7472
rect 19550 7432 19840 7460
rect 20272 7432 20536 7460
rect 20272 7401 20300 7432
rect 20530 7420 20536 7432
rect 20588 7460 20594 7472
rect 22094 7460 22100 7472
rect 20588 7432 22100 7460
rect 20588 7420 20594 7432
rect 22094 7420 22100 7432
rect 22152 7460 22158 7472
rect 23382 7460 23388 7472
rect 22152 7432 23388 7460
rect 22152 7420 22158 7432
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 21082 7352 21088 7404
rect 21140 7352 21146 7404
rect 23293 7395 23351 7401
rect 23293 7361 23305 7395
rect 23339 7392 23351 7395
rect 23842 7392 23848 7404
rect 23339 7364 23848 7392
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 18003 7296 18552 7324
rect 18003 7293 18015 7296
rect 17957 7287 18015 7293
rect 18598 7284 18604 7336
rect 18656 7324 18662 7336
rect 19981 7327 20039 7333
rect 19981 7324 19993 7327
rect 18656 7296 19993 7324
rect 18656 7284 18662 7296
rect 19981 7293 19993 7296
rect 20027 7293 20039 7327
rect 19981 7287 20039 7293
rect 21266 7284 21272 7336
rect 21324 7284 21330 7336
rect 23017 7327 23075 7333
rect 23017 7293 23029 7327
rect 23063 7324 23075 7327
rect 24854 7324 24860 7336
rect 23063 7296 24860 7324
rect 23063 7293 23075 7296
rect 23017 7287 23075 7293
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 21174 7256 21180 7268
rect 20640 7228 21180 7256
rect 20640 7188 20668 7228
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 17880 7160 20668 7188
rect 20717 7191 20775 7197
rect 17313 7151 17371 7157
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 20898 7188 20904 7200
rect 20763 7160 20904 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 18690 6984 18696 6996
rect 17460 6956 18696 6984
rect 17460 6944 17466 6956
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 13630 6916 13636 6928
rect 13412 6888 13636 6916
rect 13412 6876 13418 6888
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 16356 6888 17264 6916
rect 16356 6876 16362 6888
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6848 12587 6851
rect 12710 6848 12716 6860
rect 12575 6820 12716 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6848 12955 6851
rect 14458 6848 14464 6860
rect 12943 6820 14464 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10744 6752 10793 6780
rect 10744 6740 10750 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 11054 6672 11060 6724
rect 11112 6672 11118 6724
rect 11514 6712 11520 6724
rect 11440 6684 11520 6712
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 9766 6644 9772 6656
rect 4120 6616 9772 6644
rect 4120 6604 4126 6616
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 11440 6644 11468 6684
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 12912 6712 12940 6811
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 15988 6820 17141 6848
rect 15988 6808 15994 6820
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17236 6848 17264 6888
rect 19794 6876 19800 6928
rect 19852 6916 19858 6928
rect 20441 6919 20499 6925
rect 20441 6916 20453 6919
rect 19852 6888 20453 6916
rect 19852 6876 19858 6888
rect 20441 6885 20453 6888
rect 20487 6885 20499 6919
rect 20441 6879 20499 6885
rect 21450 6876 21456 6928
rect 21508 6916 21514 6928
rect 22830 6916 22836 6928
rect 21508 6888 22836 6916
rect 21508 6876 21514 6888
rect 22830 6876 22836 6888
rect 22888 6876 22894 6928
rect 23474 6876 23480 6928
rect 23532 6916 23538 6928
rect 23532 6888 25176 6916
rect 23532 6876 23538 6888
rect 18877 6851 18935 6857
rect 17236 6820 18644 6848
rect 17129 6811 17187 6817
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 12406 6684 12940 6712
rect 13556 6712 13584 6743
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 13780 6752 14565 6780
rect 13780 6740 13786 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 18616 6780 18644 6820
rect 18877 6817 18889 6851
rect 18923 6817 18935 6851
rect 18877 6811 18935 6817
rect 19613 6851 19671 6857
rect 19613 6817 19625 6851
rect 19659 6848 19671 6851
rect 21634 6848 21640 6860
rect 19659 6820 21640 6848
rect 19659 6817 19671 6820
rect 19613 6811 19671 6817
rect 18892 6780 18920 6811
rect 21634 6808 21640 6820
rect 21692 6808 21698 6860
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 23290 6848 23296 6860
rect 21775 6820 23296 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 25038 6808 25044 6860
rect 25096 6808 25102 6860
rect 25148 6857 25176 6888
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 21266 6780 21272 6792
rect 18616 6752 18736 6780
rect 18892 6752 21272 6780
rect 16669 6743 16727 6749
rect 14642 6712 14648 6724
rect 13556 6684 14648 6712
rect 12406 6644 12434 6684
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 14737 6715 14795 6721
rect 14737 6681 14749 6715
rect 14783 6681 14795 6715
rect 14737 6675 14795 6681
rect 15749 6715 15807 6721
rect 15749 6681 15761 6715
rect 15795 6712 15807 6715
rect 16482 6712 16488 6724
rect 15795 6684 16488 6712
rect 15795 6681 15807 6684
rect 15749 6675 15807 6681
rect 11440 6616 12434 6644
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13688 6616 13737 6644
rect 13688 6604 13694 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14366 6644 14372 6656
rect 14323 6616 14372 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14366 6604 14372 6616
rect 14424 6644 14430 6656
rect 14752 6644 14780 6675
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 14424 6616 14780 6644
rect 16684 6644 16712 6743
rect 17034 6672 17040 6724
rect 17092 6712 17098 6724
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 17092 6684 17417 6712
rect 17092 6672 17098 6684
rect 17405 6681 17417 6684
rect 17451 6712 17463 6715
rect 17678 6712 17684 6724
rect 17451 6684 17684 6712
rect 17451 6681 17463 6684
rect 17405 6675 17463 6681
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 17862 6672 17868 6724
rect 17920 6672 17926 6724
rect 18708 6712 18736 6752
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 22002 6740 22008 6792
rect 22060 6740 22066 6792
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 19797 6715 19855 6721
rect 19797 6712 19809 6715
rect 18708 6684 19809 6712
rect 19797 6681 19809 6684
rect 19843 6681 19855 6715
rect 20990 6712 20996 6724
rect 19797 6675 19855 6681
rect 20180 6684 20996 6712
rect 19150 6644 19156 6656
rect 16684 6616 19156 6644
rect 14424 6604 14430 6616
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19705 6647 19763 6653
rect 19705 6613 19717 6647
rect 19751 6644 19763 6647
rect 20070 6644 20076 6656
rect 19751 6616 20076 6644
rect 19751 6613 19763 6616
rect 19705 6607 19763 6613
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 20180 6653 20208 6684
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 21542 6672 21548 6724
rect 21600 6712 21606 6724
rect 22370 6712 22376 6724
rect 21600 6684 22376 6712
rect 21600 6672 21606 6684
rect 22370 6672 22376 6684
rect 22428 6672 22434 6724
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 24854 6712 24860 6724
rect 23891 6684 24860 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 24949 6715 25007 6721
rect 24949 6681 24961 6715
rect 24995 6712 25007 6715
rect 25222 6712 25228 6724
rect 24995 6684 25228 6712
rect 24995 6681 25007 6684
rect 24949 6675 25007 6681
rect 25222 6672 25228 6684
rect 25280 6672 25286 6724
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6613 20223 6647
rect 20165 6607 20223 6613
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 20680 6616 24593 6644
rect 20680 6604 20686 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12802 6440 12808 6452
rect 12023 6412 12808 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 14093 6443 14151 6449
rect 14093 6409 14105 6443
rect 14139 6440 14151 6443
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 14139 6412 17325 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 17313 6409 17325 6412
rect 17359 6409 17371 6443
rect 17313 6403 17371 6409
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 17920 6412 17969 6440
rect 17920 6400 17926 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 18966 6400 18972 6452
rect 19024 6440 19030 6452
rect 20622 6440 20628 6452
rect 19024 6412 20628 6440
rect 19024 6400 19030 6412
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21692 6412 22017 6440
rect 21692 6400 21698 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 23308 6412 23888 6440
rect 10689 6375 10747 6381
rect 10689 6341 10701 6375
rect 10735 6372 10747 6375
rect 11422 6372 11428 6384
rect 10735 6344 11428 6372
rect 10735 6341 10747 6344
rect 10689 6335 10747 6341
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 13872 6344 18276 6372
rect 13872 6332 13878 6344
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 6696 6276 10793 6304
rect 6696 6264 6702 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 10781 6267 10839 6273
rect 10888 6276 12081 6304
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 9364 6208 10517 6236
rect 9364 6196 9370 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 10888 6168 10916 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 12216 6276 13737 6304
rect 12216 6264 12222 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11790 6236 11796 6248
rect 11112 6208 11796 6236
rect 11112 6196 11118 6208
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 13538 6196 13544 6248
rect 13596 6196 13602 6248
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 14090 6236 14096 6248
rect 13679 6208 14096 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 14090 6196 14096 6208
rect 14148 6236 14154 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14148 6208 14381 6236
rect 14148 6196 14154 6208
rect 14369 6205 14381 6208
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16114 6236 16120 6248
rect 15887 6208 16120 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16316 6236 16344 6267
rect 17218 6264 17224 6316
rect 17276 6264 17282 6316
rect 17770 6304 17776 6316
rect 17328 6276 17776 6304
rect 17328 6236 17356 6276
rect 17770 6264 17776 6276
rect 17828 6264 17834 6316
rect 18248 6313 18276 6344
rect 19150 6332 19156 6384
rect 19208 6372 19214 6384
rect 20254 6372 20260 6384
rect 19208 6344 20260 6372
rect 19208 6332 19214 6344
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 20533 6375 20591 6381
rect 20533 6341 20545 6375
rect 20579 6372 20591 6375
rect 21542 6372 21548 6384
rect 20579 6344 21548 6372
rect 20579 6341 20591 6344
rect 20533 6335 20591 6341
rect 21542 6332 21548 6344
rect 21600 6332 21606 6384
rect 23308 6372 23336 6412
rect 23046 6344 23336 6372
rect 23382 6332 23388 6384
rect 23440 6372 23446 6384
rect 23860 6372 23888 6412
rect 24394 6400 24400 6452
rect 24452 6440 24458 6452
rect 24581 6443 24639 6449
rect 24581 6440 24593 6443
rect 24452 6412 24593 6440
rect 24452 6400 24458 6412
rect 24581 6409 24593 6412
rect 24627 6409 24639 6443
rect 24581 6403 24639 6409
rect 24670 6400 24676 6452
rect 24728 6440 24734 6452
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 24728 6412 25053 6440
rect 24728 6400 24734 6412
rect 25041 6409 25053 6412
rect 25087 6409 25099 6443
rect 25041 6403 25099 6409
rect 24688 6372 24716 6400
rect 23440 6344 23796 6372
rect 23860 6344 24716 6372
rect 23440 6332 23446 6344
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6304 19487 6307
rect 19475 6276 20668 6304
rect 19475 6273 19487 6276
rect 19429 6267 19487 6273
rect 16316 6208 17356 6236
rect 17402 6196 17408 6248
rect 17460 6196 17466 6248
rect 20640 6236 20668 6276
rect 21450 6264 21456 6316
rect 21508 6264 21514 6316
rect 23768 6313 23796 6344
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 24765 6307 24823 6313
rect 24765 6273 24777 6307
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 23382 6236 23388 6248
rect 20640 6208 23388 6236
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 23474 6196 23480 6248
rect 23532 6196 23538 6248
rect 24026 6196 24032 6248
rect 24084 6196 24090 6248
rect 6788 6140 10916 6168
rect 11149 6171 11207 6177
rect 6788 6128 6794 6140
rect 11149 6137 11161 6171
rect 11195 6168 11207 6171
rect 12526 6168 12532 6180
rect 11195 6140 12532 6168
rect 11195 6137 11207 6140
rect 11149 6131 11207 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 14550 6168 14556 6180
rect 12636 6140 14556 6168
rect 12437 6103 12495 6109
rect 12437 6069 12449 6103
rect 12483 6100 12495 6103
rect 12636 6100 12664 6140
rect 14550 6128 14556 6140
rect 14608 6128 14614 6180
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 16853 6171 16911 6177
rect 16853 6168 16865 6171
rect 14700 6140 16865 6168
rect 14700 6128 14706 6140
rect 16853 6137 16865 6140
rect 16899 6137 16911 6171
rect 24780 6168 24808 6267
rect 16853 6131 16911 6137
rect 23676 6140 24808 6168
rect 12483 6072 12664 6100
rect 12989 6103 13047 6109
rect 12483 6069 12495 6072
rect 12437 6063 12495 6069
rect 12989 6069 13001 6103
rect 13035 6100 13047 6103
rect 14458 6100 14464 6112
rect 13035 6072 14464 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 21726 6060 21732 6112
rect 21784 6100 21790 6112
rect 23676 6100 23704 6140
rect 21784 6072 23704 6100
rect 21784 6060 21790 6072
rect 24210 6060 24216 6112
rect 24268 6060 24274 6112
rect 25222 6060 25228 6112
rect 25280 6060 25286 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 11790 5856 11796 5908
rect 11848 5856 11854 5908
rect 13725 5899 13783 5905
rect 13725 5865 13737 5899
rect 13771 5896 13783 5899
rect 13814 5896 13820 5908
rect 13771 5868 13820 5896
rect 13771 5865 13783 5868
rect 13725 5859 13783 5865
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 16196 5899 16254 5905
rect 16196 5865 16208 5899
rect 16242 5896 16254 5899
rect 16850 5896 16856 5908
rect 16242 5868 16856 5896
rect 16242 5865 16254 5868
rect 16196 5859 16254 5865
rect 16850 5856 16856 5868
rect 16908 5896 16914 5908
rect 16908 5868 17264 5896
rect 16908 5856 16914 5868
rect 11422 5788 11428 5840
rect 11480 5828 11486 5840
rect 12986 5828 12992 5840
rect 11480 5800 12992 5828
rect 11480 5788 11486 5800
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13081 5831 13139 5837
rect 13081 5797 13093 5831
rect 13127 5828 13139 5831
rect 14090 5828 14096 5840
rect 13127 5800 14096 5828
rect 13127 5797 13139 5800
rect 13081 5791 13139 5797
rect 14090 5788 14096 5800
rect 14148 5788 14154 5840
rect 15473 5831 15531 5837
rect 15473 5797 15485 5831
rect 15519 5797 15531 5831
rect 17236 5828 17264 5868
rect 17678 5856 17684 5908
rect 17736 5856 17742 5908
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 17828 5868 18828 5896
rect 17828 5856 17834 5868
rect 18800 5828 18828 5868
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 23750 5896 23756 5908
rect 21508 5868 23756 5896
rect 21508 5856 21514 5868
rect 23750 5856 23756 5868
rect 23808 5856 23814 5908
rect 23845 5899 23903 5905
rect 23845 5865 23857 5899
rect 23891 5896 23903 5899
rect 24302 5896 24308 5908
rect 23891 5868 24308 5896
rect 23891 5865 23903 5868
rect 23845 5859 23903 5865
rect 24302 5856 24308 5868
rect 24360 5856 24366 5908
rect 24581 5831 24639 5837
rect 24581 5828 24593 5831
rect 17236 5800 18736 5828
rect 18800 5800 24593 5828
rect 15473 5791 15531 5797
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10778 5760 10784 5772
rect 10367 5732 10784 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 12434 5760 12440 5772
rect 11112 5732 12440 5760
rect 11112 5720 11118 5732
rect 12434 5720 12440 5732
rect 12492 5760 12498 5772
rect 14921 5763 14979 5769
rect 12492 5732 13768 5760
rect 12492 5720 12498 5732
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9640 5664 10057 5692
rect 9640 5652 9646 5664
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 11422 5652 11428 5704
rect 11480 5652 11486 5704
rect 12250 5652 12256 5704
rect 12308 5652 12314 5704
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 13446 5692 13452 5704
rect 12943 5664 13452 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 13740 5692 13768 5732
rect 14921 5729 14933 5763
rect 14967 5760 14979 5763
rect 15378 5760 15384 5772
rect 14967 5732 15384 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 15488 5760 15516 5791
rect 18708 5769 18736 5800
rect 24581 5797 24593 5800
rect 24627 5797 24639 5831
rect 24581 5791 24639 5797
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 15488 5732 18613 5760
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 19334 5720 19340 5772
rect 19392 5720 19398 5772
rect 19702 5720 19708 5772
rect 19760 5760 19766 5772
rect 24210 5760 24216 5772
rect 19760 5732 24216 5760
rect 19760 5720 19766 5732
rect 15105 5695 15163 5701
rect 15105 5692 15117 5695
rect 13740 5664 15117 5692
rect 13541 5655 13599 5661
rect 15105 5661 15117 5664
rect 15151 5661 15163 5695
rect 15105 5655 15163 5661
rect 13556 5624 13584 5655
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 19352 5692 19380 5720
rect 18555 5664 19380 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 20806 5652 20812 5704
rect 20864 5652 20870 5704
rect 22278 5652 22284 5704
rect 22336 5692 22342 5704
rect 23216 5701 23244 5732
rect 24210 5720 24216 5732
rect 24268 5720 24274 5772
rect 22465 5695 22523 5701
rect 22465 5692 22477 5695
rect 22336 5664 22477 5692
rect 22336 5652 22342 5664
rect 22465 5661 22477 5664
rect 22511 5661 22523 5695
rect 22465 5655 22523 5661
rect 23201 5695 23259 5701
rect 23201 5661 23213 5695
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 23934 5652 23940 5704
rect 23992 5692 23998 5704
rect 24029 5695 24087 5701
rect 24029 5692 24041 5695
rect 23992 5664 24041 5692
rect 23992 5652 23998 5664
rect 24029 5661 24041 5664
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 24762 5652 24768 5704
rect 24820 5652 24826 5704
rect 12452 5596 13584 5624
rect 12452 5565 12480 5596
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 14516 5596 16698 5624
rect 14516 5584 14522 5596
rect 16408 5568 16436 5596
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19613 5627 19671 5633
rect 19613 5624 19625 5627
rect 19392 5596 19625 5624
rect 19392 5584 19398 5596
rect 19613 5593 19625 5596
rect 19659 5593 19671 5627
rect 19613 5587 19671 5593
rect 20714 5584 20720 5636
rect 20772 5624 20778 5636
rect 21453 5627 21511 5633
rect 21453 5624 21465 5627
rect 20772 5596 21465 5624
rect 20772 5584 20778 5596
rect 21453 5593 21465 5596
rect 21499 5593 21511 5627
rect 21453 5587 21511 5593
rect 23385 5627 23443 5633
rect 23385 5593 23397 5627
rect 23431 5624 23443 5627
rect 23750 5624 23756 5636
rect 23431 5596 23756 5624
rect 23431 5593 23443 5596
rect 23385 5587 23443 5593
rect 23750 5584 23756 5596
rect 23808 5584 23814 5636
rect 12437 5559 12495 5565
rect 12437 5525 12449 5559
rect 12483 5525 12495 5559
rect 12437 5519 12495 5525
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 13044 5528 14289 5556
rect 13044 5516 13050 5528
rect 14277 5525 14289 5528
rect 14323 5556 14335 5559
rect 15013 5559 15071 5565
rect 15013 5556 15025 5559
rect 14323 5528 15025 5556
rect 14323 5525 14335 5528
rect 14277 5519 14335 5525
rect 15013 5525 15025 5528
rect 15059 5556 15071 5559
rect 15286 5556 15292 5568
rect 15059 5528 15292 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 16390 5516 16396 5568
rect 16448 5516 16454 5568
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5556 18199 5559
rect 18322 5556 18328 5568
rect 18187 5528 18328 5556
rect 18187 5525 18199 5528
rect 18141 5519 18199 5525
rect 18322 5516 18328 5528
rect 18380 5516 18386 5568
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 23290 5556 23296 5568
rect 22796 5528 23296 5556
rect 22796 5516 22802 5528
rect 23290 5516 23296 5528
rect 23348 5516 23354 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 22738 5352 22744 5364
rect 12636 5324 14780 5352
rect 10045 5287 10103 5293
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 11790 5284 11796 5296
rect 10091 5256 11796 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 10962 5216 10968 5228
rect 10367 5188 10968 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11146 5176 11152 5228
rect 11204 5176 11210 5228
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12636 5216 12664 5324
rect 13449 5287 13507 5293
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 13538 5284 13544 5296
rect 13495 5256 13544 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 13538 5244 13544 5256
rect 13596 5244 13602 5296
rect 14458 5244 14464 5296
rect 14516 5244 14522 5296
rect 12406 5188 12664 5216
rect 12406 5148 12434 5188
rect 12894 5176 12900 5228
rect 12952 5176 12958 5228
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 13096 5188 13185 5216
rect 10520 5120 12434 5148
rect 12529 5151 12587 5157
rect 10520 5089 10548 5120
rect 12529 5117 12541 5151
rect 12575 5148 12587 5151
rect 12912 5148 12940 5176
rect 12575 5120 12940 5148
rect 12575 5117 12587 5120
rect 12529 5111 12587 5117
rect 10505 5083 10563 5089
rect 10505 5049 10517 5083
rect 10551 5049 10563 5083
rect 10505 5043 10563 5049
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 10744 5052 12434 5080
rect 10744 5040 10750 5052
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10652 4984 10977 5012
rect 10652 4972 10658 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 12406 5012 12434 5052
rect 13096 5012 13124 5188
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 14752 5216 14780 5324
rect 18340 5324 22744 5352
rect 15286 5244 15292 5296
rect 15344 5284 15350 5296
rect 15344 5256 18000 5284
rect 15344 5244 15350 5256
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 14752 5188 15485 5216
rect 13173 5179 13231 5185
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 16942 5216 16948 5228
rect 15473 5179 15531 5185
rect 15580 5188 16948 5216
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 15580 5148 15608 5188
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 14976 5120 15608 5148
rect 14976 5108 14982 5120
rect 15746 5108 15752 5160
rect 15804 5108 15810 5160
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 17034 5148 17040 5160
rect 15896 5120 17040 5148
rect 15896 5108 15902 5120
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 17862 5108 17868 5160
rect 17920 5108 17926 5160
rect 17972 5148 18000 5256
rect 18340 5225 18368 5324
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 19794 5244 19800 5296
rect 19852 5244 19858 5296
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 20993 5287 21051 5293
rect 20993 5284 21005 5287
rect 20312 5256 21005 5284
rect 20312 5244 20318 5256
rect 20993 5253 21005 5256
rect 21039 5253 21051 5287
rect 20993 5247 21051 5253
rect 21082 5244 21088 5296
rect 21140 5284 21146 5296
rect 21140 5256 21220 5284
rect 21140 5244 21146 5256
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 20530 5176 20536 5228
rect 20588 5176 20594 5228
rect 21192 5225 21220 5256
rect 21266 5244 21272 5296
rect 21324 5284 21330 5296
rect 21545 5287 21603 5293
rect 21545 5284 21557 5287
rect 21324 5256 21557 5284
rect 21324 5244 21330 5256
rect 21545 5253 21557 5256
rect 21591 5253 21603 5287
rect 21545 5247 21603 5253
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21450 5216 21456 5228
rect 21223 5188 21456 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21450 5176 21456 5188
rect 21508 5176 21514 5228
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 23808 5188 23857 5216
rect 23808 5176 23814 5188
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 18414 5148 18420 5160
rect 17972 5120 18420 5148
rect 18414 5108 18420 5120
rect 18472 5108 18478 5160
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 18656 5120 18797 5148
rect 18656 5108 18662 5120
rect 18785 5117 18797 5120
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 20257 5151 20315 5157
rect 20257 5117 20269 5151
rect 20303 5148 20315 5151
rect 21082 5148 21088 5160
rect 20303 5120 21088 5148
rect 20303 5117 20315 5120
rect 20257 5111 20315 5117
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 21266 5108 21272 5160
rect 21324 5148 21330 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 21324 5120 22477 5148
rect 21324 5108 21330 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 23566 5108 23572 5160
rect 23624 5148 23630 5160
rect 24305 5151 24363 5157
rect 24305 5148 24317 5151
rect 23624 5120 24317 5148
rect 23624 5108 23630 5120
rect 24305 5117 24317 5120
rect 24351 5117 24363 5151
rect 24305 5111 24363 5117
rect 13906 5012 13912 5024
rect 12406 4984 13912 5012
rect 10965 4975 11023 4981
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14240 4984 14933 5012
rect 14240 4972 14246 4984
rect 14921 4981 14933 4984
rect 14967 5012 14979 5015
rect 17402 5012 17408 5024
rect 14967 4984 17408 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 22646 5012 22652 5024
rect 17736 4984 22652 5012
rect 17736 4972 17742 4984
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 14185 4811 14243 4817
rect 14185 4777 14197 4811
rect 14231 4808 14243 4811
rect 14274 4808 14280 4820
rect 14231 4780 14280 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 15212 4780 16804 4808
rect 11422 4740 11428 4752
rect 10888 4712 11428 4740
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 9582 4672 9588 4684
rect 5123 4644 9588 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 10318 4632 10324 4684
rect 10376 4632 10382 4684
rect 10594 4632 10600 4684
rect 10652 4632 10658 4684
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 1780 4576 3985 4604
rect 1780 4477 1808 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 10888 4604 10916 4712
rect 11422 4700 11428 4712
rect 11480 4700 11486 4752
rect 15212 4740 15240 4780
rect 13280 4712 15240 4740
rect 16776 4740 16804 4780
rect 16850 4768 16856 4820
rect 16908 4768 16914 4820
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 23750 4808 23756 4820
rect 17092 4780 23756 4808
rect 17092 4768 17098 4780
rect 23750 4768 23756 4780
rect 23808 4808 23814 4820
rect 24121 4811 24179 4817
rect 24121 4808 24133 4811
rect 23808 4780 24133 4808
rect 23808 4768 23814 4780
rect 24121 4777 24133 4780
rect 24167 4777 24179 4811
rect 24121 4771 24179 4777
rect 18598 4740 18604 4752
rect 16776 4712 18604 4740
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 13280 4681 13308 4712
rect 18598 4700 18604 4712
rect 18656 4700 18662 4752
rect 13265 4675 13323 4681
rect 11020 4644 12434 4672
rect 11020 4632 11026 4644
rect 7392 4576 10916 4604
rect 11057 4607 11115 4613
rect 7392 4545 7420 4576
rect 11057 4573 11069 4607
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 12406 4604 12434 4644
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 14918 4672 14924 4684
rect 13265 4635 13323 4641
rect 13372 4644 14924 4672
rect 13372 4604 13400 4644
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15105 4675 15163 4681
rect 15105 4641 15117 4675
rect 15151 4672 15163 4675
rect 15930 4672 15936 4684
rect 15151 4644 15936 4672
rect 15151 4641 15163 4644
rect 15105 4635 15163 4641
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 20530 4632 20536 4684
rect 20588 4672 20594 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 20588 4644 21281 4672
rect 20588 4632 20594 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 24581 4675 24639 4681
rect 24581 4672 24593 4675
rect 21269 4635 21327 4641
rect 22066 4644 24593 4672
rect 12406 4576 13400 4604
rect 11333 4567 11391 4573
rect 4617 4539 4675 4545
rect 4617 4505 4629 4539
rect 4663 4536 4675 4539
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 4663 4508 5365 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 6578 4508 7389 4536
rect 5353 4499 5411 4505
rect 7377 4505 7389 4508
rect 7423 4505 7435 4539
rect 7377 4499 7435 4505
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 11072 4536 11100 4567
rect 9732 4508 11100 4536
rect 11348 4536 11376 4567
rect 13722 4564 13728 4616
rect 13780 4564 13786 4616
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4604 18843 4607
rect 19610 4604 19616 4616
rect 18831 4576 19616 4604
rect 18831 4573 18843 4576
rect 18785 4567 18843 4573
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 21726 4564 21732 4616
rect 21784 4564 21790 4616
rect 21818 4564 21824 4616
rect 21876 4604 21882 4616
rect 22066 4604 22094 4644
rect 24581 4641 24593 4644
rect 24627 4641 24639 4675
rect 24581 4635 24639 4641
rect 24765 4607 24823 4613
rect 24765 4604 24777 4607
rect 21876 4576 22094 4604
rect 23584 4576 24777 4604
rect 21876 4564 21882 4576
rect 15286 4536 15292 4548
rect 11348 4508 15292 4536
rect 9732 4496 9738 4508
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 15378 4496 15384 4548
rect 15436 4496 15442 4548
rect 16390 4496 16396 4548
rect 16448 4496 16454 4548
rect 17310 4496 17316 4548
rect 17368 4536 17374 4548
rect 17589 4539 17647 4545
rect 17589 4536 17601 4539
rect 17368 4508 17601 4536
rect 17368 4496 17374 4508
rect 17589 4505 17601 4508
rect 17635 4505 17647 4539
rect 17589 4499 17647 4505
rect 20530 4496 20536 4548
rect 20588 4496 20594 4548
rect 20993 4539 21051 4545
rect 20993 4505 21005 4539
rect 21039 4536 21051 4539
rect 21634 4536 21640 4548
rect 21039 4508 21640 4536
rect 21039 4505 21051 4508
rect 20993 4499 21051 4505
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 22370 4496 22376 4548
rect 22428 4536 22434 4548
rect 22649 4539 22707 4545
rect 22649 4536 22661 4539
rect 22428 4508 22661 4536
rect 22428 4496 22434 4508
rect 22649 4505 22661 4508
rect 22695 4505 22707 4539
rect 22649 4499 22707 4505
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4437 1823 4471
rect 1765 4431 1823 4437
rect 9214 4428 9220 4480
rect 9272 4428 9278 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 11606 4468 11612 4480
rect 9539 4440 11612 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 14645 4471 14703 4477
rect 14645 4437 14657 4471
rect 14691 4468 14703 4471
rect 17218 4468 17224 4480
rect 14691 4440 17224 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 19521 4471 19579 4477
rect 19521 4437 19533 4471
rect 19567 4468 19579 4471
rect 21082 4468 21088 4480
rect 19567 4440 21088 4468
rect 19567 4437 19579 4440
rect 19521 4431 19579 4437
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 23584 4468 23612 4576
rect 24765 4573 24777 4576
rect 24811 4604 24823 4607
rect 25133 4607 25191 4613
rect 25133 4604 25145 4607
rect 24811 4576 25145 4604
rect 24811 4573 24823 4576
rect 24765 4567 24823 4573
rect 25133 4573 25145 4576
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 23750 4496 23756 4548
rect 23808 4496 23814 4548
rect 21416 4440 23612 4468
rect 21416 4428 21422 4440
rect 23658 4428 23664 4480
rect 23716 4428 23722 4480
rect 24302 4428 24308 4480
rect 24360 4468 24366 4480
rect 25317 4471 25375 4477
rect 25317 4468 25329 4471
rect 24360 4440 25329 4468
rect 24360 4428 24366 4440
rect 25317 4437 25329 4440
rect 25363 4437 25375 4471
rect 25317 4431 25375 4437
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4233 2927 4267
rect 2869 4227 2927 4233
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1544 4100 1593 4128
rect 1544 4088 1550 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 2685 4115 2743 4121
rect 2685 4081 2697 4115
rect 2731 4081 2743 4115
rect 2685 4075 2743 4081
rect 2700 3992 2728 4075
rect 2884 4060 2912 4227
rect 11146 4224 11152 4276
rect 11204 4224 11210 4276
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 15528 4236 15669 4264
rect 15528 4224 15534 4236
rect 15657 4233 15669 4236
rect 15703 4233 15715 4267
rect 15657 4227 15715 4233
rect 17862 4224 17868 4276
rect 17920 4264 17926 4276
rect 22002 4264 22008 4276
rect 17920 4236 22008 4264
rect 17920 4224 17926 4236
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 4724 4168 6040 4196
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 4120 4100 4169 4128
rect 4120 4088 4126 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4724 4128 4752 4168
rect 4157 4091 4215 4097
rect 4264 4100 4752 4128
rect 4801 4131 4859 4137
rect 4264 4060 4292 4100
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 5902 4128 5908 4140
rect 4847 4100 5908 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 6012 4128 6040 4168
rect 14182 4156 14188 4208
rect 14240 4156 14246 4208
rect 16390 4196 16396 4208
rect 15410 4168 16396 4196
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 19794 4156 19800 4208
rect 19852 4196 19858 4208
rect 20530 4196 20536 4208
rect 19852 4168 20536 4196
rect 19852 4156 19858 4168
rect 20530 4156 20536 4168
rect 20588 4196 20594 4208
rect 20588 4168 21128 4196
rect 20588 4156 20594 4168
rect 8938 4128 8944 4140
rect 6012 4100 8944 4128
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9214 4128 9220 4140
rect 9079 4100 9220 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 10226 4088 10232 4140
rect 10284 4088 10290 4140
rect 13446 4088 13452 4140
rect 13504 4088 13510 4140
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 18233 4131 18291 4137
rect 16347 4100 17264 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 7006 4060 7012 4072
rect 2884 4032 4292 4060
rect 4356 4032 7012 4060
rect 3237 3995 3295 4001
rect 3237 3992 3249 3995
rect 2700 3964 3249 3992
rect 3237 3961 3249 3964
rect 3283 3992 3295 3995
rect 3694 3992 3700 4004
rect 3283 3964 3700 3992
rect 3283 3961 3295 3964
rect 3237 3955 3295 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 4356 4001 4384 4032
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4060 11667 4063
rect 12434 4060 12440 4072
rect 11655 4032 12440 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 4341 3995 4399 4001
rect 4341 3961 4353 3995
rect 4387 3961 4399 3995
rect 4341 3955 4399 3961
rect 5353 3995 5411 4001
rect 5353 3961 5365 3995
rect 5399 3992 5411 3995
rect 5902 3992 5908 4004
rect 5399 3964 5908 3992
rect 5399 3961 5411 3964
rect 5353 3955 5411 3961
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 6604 3964 7113 3992
rect 6604 3952 6610 3964
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 10520 3992 10548 4023
rect 12434 4020 12440 4032
rect 12492 4060 12498 4072
rect 12802 4060 12808 4072
rect 12492 4032 12808 4060
rect 12492 4020 12498 4032
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 16022 4060 16028 4072
rect 13035 4032 16028 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 16264 4032 17049 4060
rect 16264 4020 16270 4032
rect 17037 4029 17049 4032
rect 17083 4029 17095 4063
rect 17236 4060 17264 4100
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18506 4128 18512 4140
rect 18279 4100 18512 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 20898 4088 20904 4140
rect 20956 4088 20962 4140
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 21100 4128 21128 4168
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 21821 4199 21879 4205
rect 21821 4196 21833 4199
rect 21508 4168 21833 4196
rect 21508 4156 21514 4168
rect 21821 4165 21833 4168
rect 21867 4165 21879 4199
rect 22097 4199 22155 4205
rect 22097 4196 22109 4199
rect 21821 4159 21879 4165
rect 21928 4168 22109 4196
rect 21637 4131 21695 4137
rect 21637 4128 21649 4131
rect 21100 4100 21649 4128
rect 21637 4097 21649 4100
rect 21683 4128 21695 4131
rect 21928 4128 21956 4168
rect 22097 4165 22109 4168
rect 22143 4196 22155 4199
rect 22465 4199 22523 4205
rect 22465 4196 22477 4199
rect 22143 4168 22477 4196
rect 22143 4165 22155 4168
rect 22097 4159 22155 4165
rect 22465 4165 22477 4168
rect 22511 4165 22523 4199
rect 22465 4159 22523 4165
rect 21683 4100 21956 4128
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 24210 4088 24216 4140
rect 24268 4088 24274 4140
rect 24302 4088 24308 4140
rect 24360 4128 24366 4140
rect 24673 4131 24731 4137
rect 24673 4128 24685 4131
rect 24360 4100 24685 4128
rect 24360 4088 24366 4100
rect 24673 4097 24685 4100
rect 24719 4097 24731 4131
rect 24673 4091 24731 4097
rect 18322 4060 18328 4072
rect 17236 4032 18328 4060
rect 17037 4023 17095 4029
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18472 4032 19165 4060
rect 18472 4020 18478 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 21082 4020 21088 4072
rect 21140 4020 21146 4072
rect 10520 3964 12434 3992
rect 7101 3955 7159 3961
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 2682 3924 2688 3936
rect 2271 3896 2688 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 3418 3884 3424 3936
rect 3476 3884 3482 3936
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4062 3924 4068 3936
rect 3927 3896 4068 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5258 3924 5264 3936
rect 5031 3896 5264 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 6089 3927 6147 3933
rect 6089 3924 6101 3927
rect 5500 3896 6101 3924
rect 5500 3884 5506 3896
rect 6089 3893 6101 3896
rect 6135 3893 6147 3927
rect 6089 3887 6147 3893
rect 7006 3884 7012 3936
rect 7064 3884 7070 3936
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7248 3896 7481 3924
rect 7248 3884 7254 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 8018 3884 8024 3936
rect 8076 3884 8082 3936
rect 9217 3927 9275 3933
rect 9217 3893 9229 3927
rect 9263 3924 9275 3927
rect 11054 3924 11060 3936
rect 9263 3896 11060 3924
rect 9263 3893 9275 3896
rect 9217 3887 9275 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 11882 3924 11888 3936
rect 11839 3896 11888 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12406 3924 12434 3964
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 16117 3995 16175 4001
rect 16117 3992 16129 3995
rect 15712 3964 16129 3992
rect 15712 3952 15718 3964
rect 16117 3961 16129 3964
rect 16163 3961 16175 3995
rect 16117 3955 16175 3961
rect 20254 3952 20260 4004
rect 20312 3992 20318 4004
rect 21266 3992 21272 4004
rect 20312 3964 21272 3992
rect 20312 3952 20318 3964
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 18874 3924 18880 3936
rect 12406 3896 18880 3924
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 20530 3884 20536 3936
rect 20588 3884 20594 3936
rect 25222 3884 25228 3936
rect 25280 3924 25286 3936
rect 25317 3927 25375 3933
rect 25317 3924 25329 3927
rect 25280 3896 25329 3924
rect 25280 3884 25286 3896
rect 25317 3893 25329 3896
rect 25363 3893 25375 3927
rect 25317 3887 25375 3893
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 1578 3680 1584 3732
rect 1636 3720 1642 3732
rect 1949 3723 2007 3729
rect 1949 3720 1961 3723
rect 1636 3692 1961 3720
rect 1636 3680 1642 3692
rect 1949 3689 1961 3692
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 7834 3720 7840 3732
rect 4479 3692 7840 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8570 3680 8576 3732
rect 8628 3680 8634 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 13814 3720 13820 3732
rect 9907 3692 13820 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 18647 3723 18705 3729
rect 18647 3689 18659 3723
rect 18693 3720 18705 3723
rect 19242 3720 19248 3732
rect 18693 3692 19248 3720
rect 18693 3689 18705 3692
rect 18647 3683 18705 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 20346 3680 20352 3732
rect 20404 3720 20410 3732
rect 22922 3720 22928 3732
rect 20404 3692 22928 3720
rect 20404 3680 20410 3692
rect 22922 3680 22928 3692
rect 22980 3680 22986 3732
rect 24029 3723 24087 3729
rect 24029 3689 24041 3723
rect 24075 3720 24087 3723
rect 24210 3720 24216 3732
rect 24075 3692 24216 3720
rect 24075 3689 24087 3692
rect 24029 3683 24087 3689
rect 24210 3680 24216 3692
rect 24268 3680 24274 3732
rect 3237 3655 3295 3661
rect 3237 3621 3249 3655
rect 3283 3652 3295 3655
rect 7466 3652 7472 3664
rect 3283 3624 7472 3652
rect 3283 3621 3295 3624
rect 3237 3615 3295 3621
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 8478 3612 8484 3664
rect 8536 3612 8542 3664
rect 10597 3655 10655 3661
rect 10597 3621 10609 3655
rect 10643 3652 10655 3655
rect 15194 3652 15200 3664
rect 10643 3624 15200 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 23382 3652 23388 3664
rect 19116 3624 23388 3652
rect 19116 3612 19122 3624
rect 23382 3612 23388 3624
rect 23440 3612 23446 3664
rect 3973 3587 4031 3593
rect 2608 3556 3648 3584
rect 2608 3525 2636 3556
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2593 3479 2651 3485
rect 2746 3488 3065 3516
rect 2222 3408 2228 3460
rect 2280 3448 2286 3460
rect 2746 3448 2774 3488
rect 3053 3485 3065 3488
rect 3099 3516 3111 3519
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3099 3488 3525 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3620 3516 3648 3556
rect 3973 3553 3985 3587
rect 4019 3584 4031 3587
rect 4798 3584 4804 3596
rect 4019 3556 4804 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 4798 3544 4804 3556
rect 4856 3584 4862 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4856 3556 4905 3584
rect 4856 3544 4862 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 8496 3584 8524 3612
rect 10870 3584 10876 3596
rect 5316 3556 8524 3584
rect 9048 3556 10876 3584
rect 5316 3544 5322 3556
rect 4154 3516 4160 3528
rect 3620 3488 4160 3516
rect 3513 3479 3571 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 6288 3488 6377 3516
rect 2280 3420 2774 3448
rect 2280 3408 2286 3420
rect 6288 3392 6316 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 7064 3488 7113 3516
rect 7064 3476 7070 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7708 3488 7757 3516
rect 7708 3476 7714 3488
rect 7745 3485 7757 3488
rect 7791 3516 7803 3519
rect 8018 3516 8024 3528
rect 7791 3488 8024 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8478 3516 8484 3528
rect 8435 3488 8484 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8478 3476 8484 3488
rect 8536 3516 8542 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8536 3488 8953 3516
rect 8536 3476 8542 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9048 3448 9076 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3584 11667 3587
rect 12066 3584 12072 3596
rect 11655 3556 12072 3584
rect 11655 3553 11667 3556
rect 11609 3547 11667 3553
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17736 3556 19901 3584
rect 17736 3544 17742 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9582 3516 9588 3528
rect 9263 3488 9588 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9582 3476 9588 3488
rect 9640 3516 9646 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9640 3488 9689 3516
rect 9640 3476 9646 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 7300 3420 9076 3448
rect 9401 3451 9459 3457
rect 1486 3340 1492 3392
rect 1544 3340 1550 3392
rect 6089 3383 6147 3389
rect 6089 3349 6101 3383
rect 6135 3380 6147 3383
rect 6270 3380 6276 3392
rect 6135 3352 6276 3380
rect 6135 3349 6147 3352
rect 6089 3343 6147 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6549 3383 6607 3389
rect 6549 3349 6561 3383
rect 6595 3380 6607 3383
rect 6638 3380 6644 3392
rect 6595 3352 6644 3380
rect 6595 3349 6607 3352
rect 6549 3343 6607 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 7300 3389 7328 3420
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 10428 3448 10456 3479
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11848 3488 11897 3516
rect 11848 3476 11854 3488
rect 11885 3485 11897 3488
rect 11931 3516 11943 3519
rect 12526 3516 12532 3528
rect 11931 3488 12532 3516
rect 11931 3485 11943 3488
rect 11885 3479 11943 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14274 3516 14280 3528
rect 13771 3488 14280 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 15654 3476 15660 3528
rect 15712 3476 15718 3528
rect 17494 3476 17500 3528
rect 17552 3476 17558 3528
rect 18874 3476 18880 3528
rect 18932 3476 18938 3528
rect 19518 3476 19524 3528
rect 19576 3476 19582 3528
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 20220 3488 21281 3516
rect 20220 3476 20226 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 21269 3479 21327 3485
rect 21836 3488 22201 3516
rect 10686 3448 10692 3460
rect 9447 3420 10692 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 12802 3408 12808 3460
rect 12860 3408 12866 3460
rect 13998 3408 14004 3460
rect 14056 3448 14062 3460
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 14056 3420 14473 3448
rect 14056 3408 14062 3420
rect 14461 3417 14473 3420
rect 14507 3417 14519 3451
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 14461 3411 14519 3417
rect 15488 3420 16313 3448
rect 15488 3392 15516 3420
rect 16301 3417 16313 3420
rect 16347 3417 16359 3451
rect 16301 3411 16359 3417
rect 18782 3408 18788 3460
rect 18840 3448 18846 3460
rect 21836 3448 21864 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 23290 3476 23296 3528
rect 23348 3516 23354 3528
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 23348 3488 23397 3516
rect 23348 3476 23354 3488
rect 23385 3485 23397 3488
rect 23431 3516 23443 3519
rect 25038 3516 25044 3528
rect 23431 3488 25044 3516
rect 23431 3485 23443 3488
rect 23385 3479 23443 3485
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 25222 3476 25228 3528
rect 25280 3476 25286 3528
rect 18840 3420 21864 3448
rect 18840 3408 18846 3420
rect 7285 3383 7343 3389
rect 7285 3349 7297 3383
rect 7331 3349 7343 3383
rect 7285 3343 7343 3349
rect 7926 3340 7932 3392
rect 7984 3340 7990 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 14734 3380 14740 3392
rect 8996 3352 14740 3380
rect 8996 3340 9002 3352
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 20990 3380 20996 3392
rect 16540 3352 20996 3380
rect 16540 3340 16546 3352
rect 20990 3340 20996 3352
rect 21048 3340 21054 3392
rect 21082 3340 21088 3392
rect 21140 3380 21146 3392
rect 22925 3383 22983 3389
rect 22925 3380 22937 3383
rect 21140 3352 22937 3380
rect 21140 3340 21146 3352
rect 22925 3349 22937 3352
rect 22971 3349 22983 3383
rect 22925 3343 22983 3349
rect 24581 3383 24639 3389
rect 24581 3349 24593 3383
rect 24627 3380 24639 3383
rect 25222 3380 25228 3392
rect 24627 3352 25228 3380
rect 24627 3349 24639 3352
rect 24581 3343 24639 3349
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4430 3176 4436 3188
rect 4304 3148 4436 3176
rect 4304 3136 4310 3148
rect 4430 3136 4436 3148
rect 4488 3176 4494 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4488 3148 4537 3176
rect 4488 3136 4494 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 6730 3136 6736 3188
rect 6788 3136 6794 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 10134 3176 10140 3188
rect 9907 3148 10140 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 15562 3176 15568 3188
rect 11195 3148 15568 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 21082 3176 21088 3188
rect 17644 3148 21088 3176
rect 17644 3136 17650 3148
rect 9401 3111 9459 3117
rect 9401 3077 9413 3111
rect 9447 3108 9459 3111
rect 11698 3108 11704 3120
rect 9447 3080 11704 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2133 3043 2191 3049
rect 2133 3040 2145 3043
rect 1903 3012 2145 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2133 3009 2145 3012
rect 2179 3040 2191 3043
rect 2590 3040 2596 3052
rect 2179 3012 2596 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3418 3000 3424 3052
rect 3476 3000 3482 3052
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 3970 3040 3976 3052
rect 3743 3012 3976 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5442 3040 5448 3052
rect 5224 3012 5448 3040
rect 5224 3000 5230 3012
rect 5442 3000 5448 3012
rect 5500 3040 5506 3052
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5500 3012 6009 3040
rect 5500 3000 5506 3012
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7800 3012 7849 3040
rect 7800 3000 7806 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8938 3040 8944 3052
rect 8159 3012 8944 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9079 3012 9689 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9677 3009 9689 3012
rect 9723 3040 9735 3043
rect 10226 3040 10232 3052
rect 9723 3012 10232 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10980 3049 11008 3080
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 15010 3108 15016 3120
rect 14292 3080 15016 3108
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 14292 3040 14320 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 20640 3117 20668 3148
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 21174 3136 21180 3188
rect 21232 3176 21238 3188
rect 21269 3179 21327 3185
rect 21269 3176 21281 3179
rect 21232 3148 21281 3176
rect 21232 3136 21238 3148
rect 21269 3145 21281 3148
rect 21315 3145 21327 3179
rect 22094 3176 22100 3188
rect 21269 3139 21327 3145
rect 22066 3136 22100 3176
rect 22152 3136 22158 3188
rect 22186 3136 22192 3188
rect 22244 3136 22250 3188
rect 22830 3136 22836 3188
rect 22888 3176 22894 3188
rect 23569 3179 23627 3185
rect 23569 3176 23581 3179
rect 22888 3148 23581 3176
rect 22888 3136 22894 3148
rect 23569 3145 23581 3148
rect 23615 3145 23627 3179
rect 23569 3139 23627 3145
rect 25038 3136 25044 3188
rect 25096 3136 25102 3188
rect 18877 3111 18935 3117
rect 18877 3108 18889 3111
rect 16632 3080 18889 3108
rect 16632 3068 16638 3080
rect 18877 3077 18889 3080
rect 18923 3077 18935 3111
rect 18877 3071 18935 3077
rect 20625 3111 20683 3117
rect 20625 3077 20637 3111
rect 20671 3077 20683 3111
rect 20625 3071 20683 3077
rect 20809 3111 20867 3117
rect 20809 3077 20821 3111
rect 20855 3108 20867 3111
rect 22066 3108 22094 3136
rect 20855 3080 22094 3108
rect 20855 3077 20867 3080
rect 20809 3071 20867 3077
rect 22738 3068 22744 3120
rect 22796 3068 22802 3120
rect 22922 3068 22928 3120
rect 22980 3108 22986 3120
rect 24213 3111 24271 3117
rect 24213 3108 24225 3111
rect 22980 3080 24225 3108
rect 22980 3068 22986 3080
rect 24213 3077 24225 3080
rect 24259 3077 24271 3111
rect 24213 3071 24271 3077
rect 24578 3068 24584 3120
rect 24636 3068 24642 3120
rect 24762 3068 24768 3120
rect 24820 3108 24826 3120
rect 25225 3111 25283 3117
rect 25225 3108 25237 3111
rect 24820 3080 25237 3108
rect 24820 3068 24826 3080
rect 25225 3077 25237 3080
rect 25271 3077 25283 3111
rect 25225 3071 25283 3077
rect 12023 3012 14320 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 1854 2904 1860 2916
rect 1719 2876 1860 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2424 2904 2452 2935
rect 5718 2932 5724 2984
rect 5776 2932 5782 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 10336 2972 10364 3003
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17184 3012 18061 3040
rect 17184 3000 17190 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 19886 3000 19892 3052
rect 19944 3000 19950 3052
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 22278 3040 22284 3052
rect 22143 3012 22284 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 22278 3000 22284 3012
rect 22336 3040 22342 3052
rect 23382 3040 23388 3052
rect 22336 3012 23388 3040
rect 22336 3000 22342 3012
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 23661 3043 23719 3049
rect 23661 3009 23673 3043
rect 23707 3040 23719 3043
rect 23707 3012 23796 3040
rect 23707 3009 23719 3012
rect 23661 3003 23719 3009
rect 11054 2972 11060 2984
rect 9263 2944 11060 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11664 2944 11713 2972
rect 11664 2932 11670 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 15896 2944 17049 2972
rect 15896 2932 15902 2944
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 21358 2932 21364 2984
rect 21416 2972 21422 2984
rect 23566 2972 23572 2984
rect 21416 2944 23572 2972
rect 21416 2932 21422 2944
rect 23566 2932 23572 2944
rect 23624 2932 23630 2984
rect 8754 2904 8760 2916
rect 2424 2876 8760 2904
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 10551 2876 12434 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 4893 2839 4951 2845
rect 4893 2805 4905 2839
rect 4939 2836 4951 2839
rect 5442 2836 5448 2848
rect 4939 2808 5448 2836
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 7377 2839 7435 2845
rect 7377 2805 7389 2839
rect 7423 2836 7435 2839
rect 11974 2836 11980 2848
rect 7423 2808 11980 2836
rect 7423 2805 7435 2808
rect 7377 2799 7435 2805
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 12406 2836 12434 2876
rect 16022 2864 16028 2916
rect 16080 2904 16086 2916
rect 23474 2904 23480 2916
rect 16080 2876 23480 2904
rect 16080 2864 16086 2876
rect 23474 2864 23480 2876
rect 23532 2864 23538 2916
rect 23768 2904 23796 3012
rect 24118 3000 24124 3052
rect 24176 3040 24182 3052
rect 25409 3043 25467 3049
rect 25409 3040 25421 3043
rect 24176 3012 25421 3040
rect 24176 3000 24182 3012
rect 25409 3009 25421 3012
rect 25455 3009 25467 3043
rect 25409 3003 25467 3009
rect 24486 2904 24492 2916
rect 23768 2876 24492 2904
rect 24486 2864 24492 2876
rect 24544 2864 24550 2916
rect 15930 2836 15936 2848
rect 12406 2808 15936 2836
rect 15930 2796 15936 2808
rect 15988 2796 15994 2848
rect 19886 2796 19892 2848
rect 19944 2836 19950 2848
rect 22370 2836 22376 2848
rect 19944 2808 22376 2836
rect 19944 2796 19950 2808
rect 22370 2796 22376 2808
rect 22428 2796 22434 2848
rect 23382 2796 23388 2848
rect 23440 2836 23446 2848
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23440 2808 24133 2836
rect 23440 2796 23446 2808
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 24121 2799 24179 2805
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4617 2635 4675 2641
rect 4617 2632 4629 2635
rect 4212 2604 4629 2632
rect 4212 2592 4218 2604
rect 4617 2601 4629 2604
rect 4663 2601 4675 2635
rect 4617 2595 4675 2601
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 9122 2632 9128 2644
rect 6871 2604 9128 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 13906 2632 13912 2644
rect 9355 2604 13912 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 14366 2632 14372 2644
rect 14231 2604 14372 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 16393 2635 16451 2641
rect 16393 2632 16405 2635
rect 16255 2604 16405 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 16393 2601 16405 2604
rect 16439 2632 16451 2635
rect 16482 2632 16488 2644
rect 16439 2604 16488 2632
rect 16439 2601 16451 2604
rect 16393 2595 16451 2601
rect 16482 2592 16488 2604
rect 16540 2592 16546 2644
rect 18693 2635 18751 2641
rect 18693 2601 18705 2635
rect 18739 2632 18751 2635
rect 18874 2632 18880 2644
rect 18739 2604 18880 2632
rect 18739 2601 18751 2604
rect 18693 2595 18751 2601
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 23198 2632 23204 2644
rect 20496 2604 23204 2632
rect 20496 2592 20502 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 23845 2635 23903 2641
rect 23845 2632 23857 2635
rect 23716 2604 23857 2632
rect 23716 2592 23722 2604
rect 23845 2601 23857 2604
rect 23891 2601 23903 2635
rect 23845 2595 23903 2601
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 9674 2564 9680 2576
rect 7975 2536 9680 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 12158 2564 12164 2576
rect 9784 2536 12164 2564
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 2832 2468 4016 2496
rect 2832 2456 2838 2468
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 1854 2428 1860 2440
rect 1719 2400 1860 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2363 2400 2605 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2593 2397 2605 2400
rect 2639 2428 2651 2431
rect 2639 2400 2774 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2746 2360 2774 2400
rect 2866 2388 2872 2440
rect 2924 2388 2930 2440
rect 3988 2437 4016 2468
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5316 2468 5457 2496
rect 5316 2456 5322 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 8846 2496 8852 2508
rect 5445 2459 5503 2465
rect 7116 2468 8852 2496
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5350 2428 5356 2440
rect 5215 2400 5356 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 7116 2437 7144 2468
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 9784 2496 9812 2536
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 15746 2564 15752 2576
rect 12406 2536 15752 2564
rect 9048 2468 9812 2496
rect 10689 2499 10747 2505
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6503 2400 7113 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 8294 2428 8300 2440
rect 7791 2400 8300 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 9048 2428 9076 2468
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 10962 2496 10968 2508
rect 10735 2468 10968 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 12406 2496 12434 2536
rect 15746 2524 15752 2536
rect 15804 2524 15810 2576
rect 16114 2524 16120 2576
rect 16172 2564 16178 2576
rect 22186 2564 22192 2576
rect 16172 2536 22192 2564
rect 16172 2524 16178 2536
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 11164 2468 12434 2496
rect 8389 2391 8447 2397
rect 8496 2400 9076 2428
rect 2958 2360 2964 2372
rect 2746 2332 2964 2360
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 7834 2360 7840 2372
rect 6687 2332 7840 2360
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 7834 2320 7840 2332
rect 7892 2360 7898 2372
rect 8404 2360 8432 2391
rect 7892 2332 8432 2360
rect 7892 2320 7898 2332
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 7098 2292 7104 2304
rect 1903 2264 7104 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7285 2295 7343 2301
rect 7285 2261 7297 2295
rect 7331 2292 7343 2295
rect 8496 2292 8524 2400
rect 9122 2388 9128 2440
rect 9180 2428 9186 2440
rect 9950 2428 9956 2440
rect 9180 2400 9956 2428
rect 9180 2388 9186 2400
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 11164 2437 11192 2468
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15160 2468 17325 2496
rect 15160 2456 15166 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 17313 2459 17371 2465
rect 17972 2468 19901 2496
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2428 11759 2431
rect 11882 2428 11888 2440
rect 11747 2400 11888 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14148 2400 14473 2428
rect 14148 2388 14154 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17972 2428 18000 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 20956 2468 21281 2496
rect 20956 2456 20962 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 24762 2496 24768 2508
rect 21269 2459 21327 2465
rect 23400 2468 24768 2496
rect 17000 2400 18000 2428
rect 18877 2431 18935 2437
rect 17000 2388 17006 2400
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19058 2428 19064 2440
rect 18923 2400 19064 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19518 2388 19524 2440
rect 19576 2428 19582 2440
rect 23400 2437 23428 2468
rect 24762 2456 24768 2468
rect 24820 2456 24826 2508
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 19576 2400 22201 2428
rect 19576 2388 19582 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2428 24087 2431
rect 24118 2428 24124 2440
rect 24075 2400 24124 2428
rect 24075 2397 24087 2400
rect 24029 2391 24087 2397
rect 24118 2388 24124 2400
rect 24176 2388 24182 2440
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 12342 2360 12348 2372
rect 8588 2332 12348 2360
rect 8588 2301 8616 2332
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 16298 2360 16304 2372
rect 16040 2332 16304 2360
rect 7331 2264 8524 2292
rect 8573 2295 8631 2301
rect 7331 2261 7343 2264
rect 7285 2255 7343 2261
rect 8573 2261 8585 2295
rect 8619 2261 8631 2295
rect 8573 2255 8631 2261
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 16040 2292 16068 2332
rect 16298 2320 16304 2332
rect 16356 2320 16362 2372
rect 11931 2264 16068 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 24578 2252 24584 2304
rect 24636 2252 24642 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 9766 2088 9772 2100
rect 2924 2060 9772 2088
rect 2924 2048 2930 2060
rect 9766 2048 9772 2060
rect 9824 2048 9830 2100
rect 8294 1980 8300 2032
rect 8352 2020 8358 2032
rect 20530 2020 20536 2032
rect 8352 1992 20536 2020
rect 8352 1980 8358 1992
rect 20530 1980 20536 1992
rect 20588 1980 20594 2032
rect 7650 1912 7656 1964
rect 7708 1952 7714 1964
rect 24578 1952 24584 1964
rect 7708 1924 24584 1952
rect 7708 1912 7714 1924
rect 24578 1912 24584 1924
rect 24636 1912 24642 1964
rect 10962 1844 10968 1896
rect 11020 1884 11026 1896
rect 22094 1884 22100 1896
rect 11020 1856 22100 1884
rect 11020 1844 11026 1856
rect 22094 1844 22100 1856
rect 22152 1844 22158 1896
rect 7098 1776 7104 1828
rect 7156 1816 7162 1828
rect 11330 1816 11336 1828
rect 7156 1788 11336 1816
rect 7156 1776 7162 1788
rect 11330 1776 11336 1788
rect 11388 1776 11394 1828
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 13820 54315 13872 54324
rect 13820 54281 13829 54315
rect 13829 54281 13863 54315
rect 13863 54281 13872 54315
rect 13820 54272 13872 54281
rect 18972 54315 19024 54324
rect 18972 54281 18981 54315
rect 18981 54281 19015 54315
rect 19015 54281 19024 54315
rect 18972 54272 19024 54281
rect 2412 54247 2464 54256
rect 2412 54213 2421 54247
rect 2421 54213 2455 54247
rect 2455 54213 2464 54247
rect 2412 54204 2464 54213
rect 5172 54204 5224 54256
rect 4988 54136 5040 54188
rect 6000 54179 6052 54188
rect 6000 54145 6009 54179
rect 6009 54145 6043 54179
rect 6043 54145 6052 54179
rect 6000 54136 6052 54145
rect 8392 54179 8444 54188
rect 8392 54145 8401 54179
rect 8401 54145 8435 54179
rect 8435 54145 8444 54179
rect 8392 54136 8444 54145
rect 9588 54179 9640 54188
rect 9588 54145 9597 54179
rect 9597 54145 9631 54179
rect 9631 54145 9640 54179
rect 9588 54136 9640 54145
rect 11704 54136 11756 54188
rect 7840 54111 7892 54120
rect 7840 54077 7849 54111
rect 7849 54077 7883 54111
rect 7883 54077 7892 54111
rect 7840 54068 7892 54077
rect 9312 54068 9364 54120
rect 12348 54068 12400 54120
rect 14832 54136 14884 54188
rect 16580 54136 16632 54188
rect 17592 54136 17644 54188
rect 20720 54136 20772 54188
rect 22100 54136 22152 54188
rect 8484 54000 8536 54052
rect 25872 54136 25924 54188
rect 13912 54000 13964 54052
rect 16764 54000 16816 54052
rect 12716 53932 12768 53984
rect 16856 53975 16908 53984
rect 16856 53941 16865 53975
rect 16865 53941 16899 53975
rect 16899 53941 16908 53975
rect 16856 53932 16908 53941
rect 17500 53932 17552 53984
rect 22100 53975 22152 53984
rect 22100 53941 22109 53975
rect 22109 53941 22143 53975
rect 22143 53941 22152 53975
rect 22100 53932 22152 53941
rect 24676 53932 24728 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 10692 53660 10744 53712
rect 1032 53592 1084 53644
rect 3792 53592 3844 53644
rect 6552 53592 6604 53644
rect 24860 53660 24912 53712
rect 23296 53592 23348 53644
rect 5356 53567 5408 53576
rect 5356 53533 5365 53567
rect 5365 53533 5399 53567
rect 5399 53533 5408 53567
rect 5356 53524 5408 53533
rect 9220 53524 9272 53576
rect 10692 53524 10744 53576
rect 22560 53567 22612 53576
rect 22560 53533 22569 53567
rect 22569 53533 22603 53567
rect 22603 53533 22612 53567
rect 22560 53524 22612 53533
rect 23388 53524 23440 53576
rect 24676 53567 24728 53576
rect 24676 53533 24685 53567
rect 24685 53533 24719 53567
rect 24719 53533 24728 53567
rect 24676 53524 24728 53533
rect 5540 53456 5592 53508
rect 22744 53456 22796 53508
rect 22652 53388 22704 53440
rect 23664 53388 23716 53440
rect 24584 53388 24636 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 4988 53184 5040 53236
rect 22560 53184 22612 53236
rect 23296 53227 23348 53236
rect 23296 53193 23305 53227
rect 23305 53193 23339 53227
rect 23339 53193 23348 53227
rect 23296 53184 23348 53193
rect 23388 53227 23440 53236
rect 23388 53193 23397 53227
rect 23397 53193 23431 53227
rect 23431 53193 23440 53227
rect 23388 53184 23440 53193
rect 24768 53184 24820 53236
rect 25320 53227 25372 53236
rect 25320 53193 25329 53227
rect 25329 53193 25363 53227
rect 25363 53193 25372 53227
rect 25320 53184 25372 53193
rect 7564 53048 7616 53100
rect 25504 52955 25556 52964
rect 25504 52921 25513 52955
rect 25513 52921 25547 52955
rect 25547 52921 25556 52955
rect 25504 52912 25556 52921
rect 23848 52887 23900 52896
rect 23848 52853 23857 52887
rect 23857 52853 23891 52887
rect 23891 52853 23900 52887
rect 23848 52844 23900 52853
rect 24124 52844 24176 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 5356 52640 5408 52692
rect 24492 52683 24544 52692
rect 24492 52649 24501 52683
rect 24501 52649 24535 52683
rect 24535 52649 24544 52683
rect 24492 52640 24544 52649
rect 23572 52572 23624 52624
rect 17408 52504 17460 52556
rect 9404 52436 9456 52488
rect 24492 52436 24544 52488
rect 25228 52411 25280 52420
rect 25228 52377 25237 52411
rect 25237 52377 25271 52411
rect 25271 52377 25280 52411
rect 25228 52368 25280 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 25228 52096 25280 52148
rect 24584 52003 24636 52012
rect 24584 51969 24593 52003
rect 24593 51969 24627 52003
rect 24627 51969 24636 52003
rect 24584 51960 24636 51969
rect 25504 51960 25556 52012
rect 24400 51799 24452 51808
rect 24400 51765 24409 51799
rect 24409 51765 24443 51799
rect 24443 51765 24452 51799
rect 24400 51756 24452 51765
rect 26884 51756 26936 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 8392 51552 8444 51604
rect 9220 51595 9272 51604
rect 9220 51561 9229 51595
rect 9229 51561 9263 51595
rect 9263 51561 9272 51595
rect 9220 51552 9272 51561
rect 6000 51484 6052 51536
rect 7840 51348 7892 51400
rect 10416 51348 10468 51400
rect 10324 51280 10376 51332
rect 25228 51323 25280 51332
rect 25228 51289 25237 51323
rect 25237 51289 25271 51323
rect 25271 51289 25280 51323
rect 25228 51280 25280 51289
rect 26516 51212 26568 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 25228 50915 25280 50924
rect 25228 50881 25237 50915
rect 25237 50881 25271 50915
rect 25271 50881 25280 50915
rect 25228 50872 25280 50881
rect 26240 50668 26292 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 5540 50464 5592 50516
rect 6644 50464 6696 50516
rect 8484 50464 8536 50516
rect 9588 50507 9640 50516
rect 9588 50473 9597 50507
rect 9597 50473 9631 50507
rect 9631 50473 9640 50507
rect 9588 50464 9640 50473
rect 7564 50439 7616 50448
rect 7564 50405 7573 50439
rect 7573 50405 7607 50439
rect 7607 50405 7616 50439
rect 7564 50396 7616 50405
rect 9496 50396 9548 50448
rect 8484 50260 8536 50312
rect 9588 50260 9640 50312
rect 25320 50124 25372 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 25136 49716 25188 49768
rect 25320 49759 25372 49768
rect 25320 49725 25329 49759
rect 25329 49725 25363 49759
rect 25363 49725 25372 49759
rect 25320 49716 25372 49725
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 10692 49351 10744 49360
rect 10692 49317 10701 49351
rect 10701 49317 10735 49351
rect 10735 49317 10744 49351
rect 10692 49308 10744 49317
rect 11704 49351 11756 49360
rect 11704 49317 11713 49351
rect 11713 49317 11747 49351
rect 11747 49317 11756 49351
rect 11704 49308 11756 49317
rect 10232 49104 10284 49156
rect 10968 49104 11020 49156
rect 25228 49147 25280 49156
rect 25228 49113 25237 49147
rect 25237 49113 25271 49147
rect 25271 49113 25280 49147
rect 25228 49104 25280 49113
rect 25596 49036 25648 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 6644 48875 6696 48884
rect 6644 48841 6653 48875
rect 6653 48841 6687 48875
rect 6687 48841 6696 48875
rect 6644 48832 6696 48841
rect 8668 48764 8720 48816
rect 8852 48560 8904 48612
rect 8668 48535 8720 48544
rect 8668 48501 8677 48535
rect 8677 48501 8711 48535
rect 8711 48501 8720 48535
rect 8668 48492 8720 48501
rect 10876 48492 10928 48544
rect 25228 48492 25280 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 9496 48084 9548 48136
rect 24400 48084 24452 48136
rect 25228 48127 25280 48136
rect 25228 48093 25237 48127
rect 25237 48093 25271 48127
rect 25271 48093 25280 48127
rect 25228 48084 25280 48093
rect 12624 47948 12676 48000
rect 21824 47948 21876 48000
rect 25872 47948 25924 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9404 47744 9456 47796
rect 8484 47676 8536 47728
rect 10784 47676 10836 47728
rect 25320 47651 25372 47660
rect 25320 47617 25329 47651
rect 25329 47617 25363 47651
rect 25363 47617 25372 47651
rect 25320 47608 25372 47617
rect 8852 47404 8904 47456
rect 9128 47404 9180 47456
rect 25412 47404 25464 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 9404 46996 9456 47048
rect 13728 46928 13780 46980
rect 25320 46860 25372 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 9772 46656 9824 46708
rect 10324 46699 10376 46708
rect 10324 46665 10333 46699
rect 10333 46665 10367 46699
rect 10367 46665 10376 46699
rect 10324 46656 10376 46665
rect 10784 46656 10836 46708
rect 11060 46699 11112 46708
rect 11060 46665 11069 46699
rect 11069 46665 11103 46699
rect 11103 46665 11112 46699
rect 11060 46656 11112 46665
rect 10784 46563 10836 46572
rect 10784 46529 10793 46563
rect 10793 46529 10827 46563
rect 10827 46529 10836 46563
rect 10784 46520 10836 46529
rect 13728 46588 13780 46640
rect 13912 46563 13964 46572
rect 13912 46529 13921 46563
rect 13921 46529 13955 46563
rect 13955 46529 13964 46563
rect 13912 46520 13964 46529
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 15752 46495 15804 46504
rect 15752 46461 15761 46495
rect 15761 46461 15795 46495
rect 15795 46461 15804 46495
rect 15752 46452 15804 46461
rect 10600 46359 10652 46368
rect 10600 46325 10609 46359
rect 10609 46325 10643 46359
rect 10643 46325 10652 46359
rect 10600 46316 10652 46325
rect 16488 46316 16540 46368
rect 25044 46316 25096 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 7840 46112 7892 46164
rect 9496 45976 9548 46028
rect 21732 46044 21784 46096
rect 16856 45976 16908 46028
rect 8576 45951 8628 45960
rect 8576 45917 8585 45951
rect 8585 45917 8619 45951
rect 8619 45917 8628 45951
rect 8576 45908 8628 45917
rect 10416 45908 10468 45960
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 16488 45883 16540 45892
rect 16488 45849 16497 45883
rect 16497 45849 16531 45883
rect 16531 45849 16540 45883
rect 16488 45840 16540 45849
rect 15108 45772 15160 45824
rect 24952 45772 25004 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 12624 45500 12676 45552
rect 12716 45475 12768 45484
rect 12716 45441 12725 45475
rect 12725 45441 12759 45475
rect 12759 45441 12768 45475
rect 12716 45432 12768 45441
rect 14556 45407 14608 45416
rect 14556 45373 14565 45407
rect 14565 45373 14599 45407
rect 14599 45373 14608 45407
rect 14556 45364 14608 45373
rect 25320 45228 25372 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 9128 45067 9180 45076
rect 9128 45033 9137 45067
rect 9137 45033 9171 45067
rect 9171 45033 9180 45067
rect 9128 45024 9180 45033
rect 19984 44956 20036 45008
rect 17500 44931 17552 44940
rect 17500 44897 17509 44931
rect 17509 44897 17543 44931
rect 17543 44897 17552 44931
rect 17500 44888 17552 44897
rect 10876 44863 10928 44872
rect 10876 44829 10885 44863
rect 10885 44829 10919 44863
rect 10919 44829 10928 44863
rect 10876 44820 10928 44829
rect 8668 44684 8720 44736
rect 10600 44795 10652 44804
rect 10600 44761 10609 44795
rect 10609 44761 10643 44795
rect 10643 44761 10652 44795
rect 10600 44752 10652 44761
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 15108 44752 15160 44804
rect 11152 44727 11204 44736
rect 11152 44693 11161 44727
rect 11161 44693 11195 44727
rect 11195 44693 11204 44727
rect 11152 44684 11204 44693
rect 11336 44727 11388 44736
rect 11336 44693 11345 44727
rect 11345 44693 11379 44727
rect 11379 44693 11388 44727
rect 11336 44684 11388 44693
rect 25320 44684 25372 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 9588 44523 9640 44532
rect 9588 44489 9597 44523
rect 9597 44489 9631 44523
rect 9631 44489 9640 44523
rect 9588 44480 9640 44489
rect 9220 44344 9272 44396
rect 11060 44387 11112 44396
rect 11060 44353 11069 44387
rect 11069 44353 11103 44387
rect 11103 44353 11112 44387
rect 11060 44344 11112 44353
rect 25228 44387 25280 44396
rect 25228 44353 25237 44387
rect 25237 44353 25271 44387
rect 25271 44353 25280 44387
rect 25228 44344 25280 44353
rect 8944 44319 8996 44328
rect 8944 44285 8953 44319
rect 8953 44285 8987 44319
rect 8987 44285 8996 44319
rect 8944 44276 8996 44285
rect 10416 44140 10468 44192
rect 10968 44183 11020 44192
rect 10968 44149 10977 44183
rect 10977 44149 11011 44183
rect 11011 44149 11020 44183
rect 10968 44140 11020 44149
rect 25688 44140 25740 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 21824 43843 21876 43852
rect 21824 43809 21833 43843
rect 21833 43809 21867 43843
rect 21867 43809 21876 43843
rect 21824 43800 21876 43809
rect 20720 43732 20772 43784
rect 23388 43732 23440 43784
rect 16580 43596 16632 43648
rect 25228 43596 25280 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 25228 43299 25280 43308
rect 25228 43265 25237 43299
rect 25237 43265 25271 43299
rect 25271 43265 25280 43299
rect 25228 43256 25280 43265
rect 24308 43120 24360 43172
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 9772 42755 9824 42764
rect 9772 42721 9781 42755
rect 9781 42721 9815 42755
rect 9815 42721 9824 42755
rect 9772 42712 9824 42721
rect 10232 42755 10284 42764
rect 10232 42721 10241 42755
rect 10241 42721 10275 42755
rect 10275 42721 10284 42755
rect 10232 42712 10284 42721
rect 9036 42644 9088 42696
rect 25228 42619 25280 42628
rect 25228 42585 25237 42619
rect 25237 42585 25271 42619
rect 25271 42585 25280 42619
rect 25228 42576 25280 42585
rect 20996 42508 21048 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 10600 42304 10652 42356
rect 11152 42304 11204 42356
rect 11520 42304 11572 42356
rect 10968 42236 11020 42288
rect 11336 42100 11388 42152
rect 11520 42007 11572 42016
rect 11520 41973 11529 42007
rect 11529 41973 11563 42007
rect 11563 41973 11572 42007
rect 11520 41964 11572 41973
rect 11704 42007 11756 42016
rect 11704 41973 11713 42007
rect 11713 41973 11747 42007
rect 11747 41973 11756 42007
rect 11704 41964 11756 41973
rect 25228 41964 25280 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 10876 41803 10928 41812
rect 10876 41769 10885 41803
rect 10885 41769 10919 41803
rect 10919 41769 10928 41803
rect 10876 41760 10928 41769
rect 10416 41667 10468 41676
rect 10416 41633 10425 41667
rect 10425 41633 10459 41667
rect 10459 41633 10468 41667
rect 10416 41624 10468 41633
rect 10232 41599 10284 41608
rect 10232 41565 10241 41599
rect 10241 41565 10275 41599
rect 10275 41565 10284 41599
rect 10232 41556 10284 41565
rect 25228 41599 25280 41608
rect 25228 41565 25237 41599
rect 25237 41565 25271 41599
rect 25271 41565 25280 41599
rect 25228 41556 25280 41565
rect 24860 41488 24912 41540
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 24860 40876 24912 40928
rect 25044 40876 25096 40928
rect 26608 40876 26660 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 24952 40332 25004 40384
rect 25228 40332 25280 40384
rect 25504 40375 25556 40384
rect 25504 40341 25513 40375
rect 25513 40341 25547 40375
rect 25547 40341 25556 40375
rect 25504 40332 25556 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 23296 40128 23348 40180
rect 25504 40060 25556 40112
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 22008 39244 22060 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 25320 38700 25372 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 25320 38335 25372 38344
rect 25320 38301 25329 38335
rect 25329 38301 25363 38335
rect 25363 38301 25372 38335
rect 25320 38292 25372 38301
rect 25504 38156 25556 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 8576 37952 8628 38004
rect 8852 37859 8904 37868
rect 8852 37825 8861 37859
rect 8861 37825 8895 37859
rect 8895 37825 8904 37859
rect 8852 37816 8904 37825
rect 25228 37859 25280 37868
rect 25228 37825 25237 37859
rect 25237 37825 25271 37859
rect 25271 37825 25280 37859
rect 25228 37816 25280 37825
rect 25964 37612 26016 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 25228 37068 25280 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 25228 36771 25280 36780
rect 25228 36737 25237 36771
rect 25237 36737 25271 36771
rect 25271 36737 25280 36771
rect 25228 36728 25280 36737
rect 25780 36524 25832 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 26792 35980 26844 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 11704 35776 11756 35828
rect 25044 35776 25096 35828
rect 11520 35751 11572 35760
rect 11520 35717 11529 35751
rect 11529 35717 11563 35751
rect 11563 35717 11572 35751
rect 11520 35708 11572 35717
rect 24860 35708 24912 35760
rect 15752 35640 15804 35692
rect 21088 35683 21140 35692
rect 21088 35649 21097 35683
rect 21097 35649 21131 35683
rect 21131 35649 21140 35683
rect 21088 35640 21140 35649
rect 21732 35640 21784 35692
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 10968 35572 11020 35624
rect 21272 35615 21324 35624
rect 21272 35581 21281 35615
rect 21281 35581 21315 35615
rect 21315 35581 21324 35615
rect 21272 35572 21324 35581
rect 22560 35615 22612 35624
rect 22560 35581 22569 35615
rect 22569 35581 22603 35615
rect 22603 35581 22612 35615
rect 22560 35572 22612 35581
rect 19248 35504 19300 35556
rect 11796 35479 11848 35488
rect 11796 35445 11805 35479
rect 11805 35445 11839 35479
rect 11839 35445 11848 35479
rect 11796 35436 11848 35445
rect 20536 35504 20588 35556
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 21732 35232 21784 35284
rect 22284 35096 22336 35148
rect 24952 35028 25004 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 19984 34960 20036 35012
rect 20260 34960 20312 35012
rect 22744 34935 22796 34944
rect 22744 34901 22753 34935
rect 22753 34901 22787 34935
rect 22787 34901 22796 34935
rect 22744 34892 22796 34901
rect 26148 34892 26200 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 20352 34688 20404 34740
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 20720 34348 20772 34400
rect 21824 34348 21876 34400
rect 22192 34348 22244 34400
rect 22652 34348 22704 34400
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 8944 34144 8996 34196
rect 22100 34144 22152 34196
rect 22560 34144 22612 34196
rect 11796 34008 11848 34060
rect 22652 34008 22704 34060
rect 23388 34051 23440 34060
rect 23388 34017 23397 34051
rect 23397 34017 23431 34051
rect 23431 34017 23440 34051
rect 23388 34008 23440 34017
rect 9220 33940 9272 33992
rect 19340 33940 19392 33992
rect 16304 33872 16356 33924
rect 19708 33915 19760 33924
rect 19708 33881 19717 33915
rect 19717 33881 19751 33915
rect 19751 33881 19760 33915
rect 19708 33872 19760 33881
rect 20168 33872 20220 33924
rect 21824 33872 21876 33924
rect 23204 33872 23256 33924
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 21180 33847 21232 33856
rect 21180 33813 21189 33847
rect 21189 33813 21223 33847
rect 21223 33813 21232 33847
rect 21180 33804 21232 33813
rect 24216 33804 24268 33856
rect 26240 33804 26292 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 20168 33600 20220 33652
rect 21824 33600 21876 33652
rect 22284 33575 22336 33584
rect 22284 33541 22293 33575
rect 22293 33541 22327 33575
rect 22327 33541 22336 33575
rect 22284 33532 22336 33541
rect 22560 33600 22612 33652
rect 19708 33260 19760 33312
rect 20444 33260 20496 33312
rect 23296 33396 23348 33448
rect 22100 33260 22152 33312
rect 24216 33303 24268 33312
rect 24216 33269 24225 33303
rect 24225 33269 24259 33303
rect 24259 33269 24268 33303
rect 24216 33260 24268 33269
rect 24584 33303 24636 33312
rect 24584 33269 24593 33303
rect 24593 33269 24627 33303
rect 24627 33269 24636 33303
rect 24584 33260 24636 33269
rect 24768 33260 24820 33312
rect 25412 33328 25464 33380
rect 26424 33328 26476 33380
rect 26056 33260 26108 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 16764 33099 16816 33108
rect 16764 33065 16773 33099
rect 16773 33065 16807 33099
rect 16807 33065 16816 33099
rect 16764 33056 16816 33065
rect 17316 33056 17368 33108
rect 22284 33099 22336 33108
rect 22284 33065 22293 33099
rect 22293 33065 22327 33099
rect 22327 33065 22336 33099
rect 22284 33056 22336 33065
rect 23572 33056 23624 33108
rect 16212 32963 16264 32972
rect 16212 32929 16221 32963
rect 16221 32929 16255 32963
rect 16255 32929 16264 32963
rect 16580 32963 16632 32972
rect 16212 32920 16264 32929
rect 16580 32929 16589 32963
rect 16589 32929 16623 32963
rect 16623 32929 16632 32963
rect 16580 32920 16632 32929
rect 16764 32852 16816 32904
rect 12624 32716 12676 32768
rect 23296 32920 23348 32972
rect 24952 32920 25004 32972
rect 26608 32852 26660 32904
rect 17224 32716 17276 32768
rect 20812 32784 20864 32836
rect 23204 32784 23256 32836
rect 25412 32784 25464 32836
rect 21824 32716 21876 32768
rect 24584 32716 24636 32768
rect 25228 32716 25280 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 16672 32512 16724 32564
rect 23848 32512 23900 32564
rect 16304 32487 16356 32496
rect 16304 32453 16313 32487
rect 16313 32453 16347 32487
rect 16347 32453 16356 32487
rect 16304 32444 16356 32453
rect 20076 32444 20128 32496
rect 21180 32444 21232 32496
rect 23204 32444 23256 32496
rect 23756 32444 23808 32496
rect 24216 32444 24268 32496
rect 15476 32351 15528 32360
rect 15476 32317 15485 32351
rect 15485 32317 15519 32351
rect 15519 32317 15528 32351
rect 15476 32308 15528 32317
rect 21824 32376 21876 32428
rect 22468 32376 22520 32428
rect 23296 32376 23348 32428
rect 20812 32351 20864 32360
rect 17040 32215 17092 32224
rect 17040 32181 17049 32215
rect 17049 32181 17083 32215
rect 17083 32181 17092 32215
rect 17040 32172 17092 32181
rect 19064 32215 19116 32224
rect 19064 32181 19073 32215
rect 19073 32181 19107 32215
rect 19107 32181 19116 32215
rect 19064 32172 19116 32181
rect 19432 32172 19484 32224
rect 20812 32317 20821 32351
rect 20821 32317 20855 32351
rect 20855 32317 20864 32351
rect 20812 32308 20864 32317
rect 24952 32308 25004 32360
rect 21088 32215 21140 32224
rect 21088 32181 21097 32215
rect 21097 32181 21131 32215
rect 21131 32181 21140 32215
rect 21088 32172 21140 32181
rect 21824 32172 21876 32224
rect 22100 32172 22152 32224
rect 22836 32172 22888 32224
rect 25412 32172 25464 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 16856 31968 16908 32020
rect 17408 31968 17460 32020
rect 20168 31968 20220 32020
rect 21088 31968 21140 32020
rect 12532 31900 12584 31952
rect 16212 31875 16264 31884
rect 16212 31841 16221 31875
rect 16221 31841 16255 31875
rect 16255 31841 16264 31875
rect 16212 31832 16264 31841
rect 17776 31832 17828 31884
rect 19708 31875 19760 31884
rect 19708 31841 19717 31875
rect 19717 31841 19751 31875
rect 19751 31841 19760 31875
rect 19708 31832 19760 31841
rect 20904 31832 20956 31884
rect 22008 31832 22060 31884
rect 22836 31900 22888 31952
rect 25044 31900 25096 31952
rect 23388 31832 23440 31884
rect 15476 31764 15528 31816
rect 16764 31807 16816 31816
rect 16764 31773 16773 31807
rect 16773 31773 16807 31807
rect 16807 31773 16816 31807
rect 16764 31764 16816 31773
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 23020 31764 23072 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 17132 31696 17184 31748
rect 20168 31696 20220 31748
rect 16672 31628 16724 31680
rect 18788 31671 18840 31680
rect 18788 31637 18797 31671
rect 18797 31637 18831 31671
rect 18831 31637 18840 31671
rect 18788 31628 18840 31637
rect 21640 31671 21692 31680
rect 21640 31637 21649 31671
rect 21649 31637 21683 31671
rect 21683 31637 21692 31671
rect 21640 31628 21692 31637
rect 22008 31671 22060 31680
rect 22008 31637 22017 31671
rect 22017 31637 22051 31671
rect 22051 31637 22060 31671
rect 22008 31628 22060 31637
rect 22376 31628 22428 31680
rect 22652 31671 22704 31680
rect 22652 31637 22661 31671
rect 22661 31637 22695 31671
rect 22695 31637 22704 31671
rect 22652 31628 22704 31637
rect 24032 31671 24084 31680
rect 24032 31637 24041 31671
rect 24041 31637 24075 31671
rect 24075 31637 24084 31671
rect 24032 31628 24084 31637
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 14464 31356 14516 31408
rect 16212 31424 16264 31476
rect 17132 31424 17184 31476
rect 16764 31288 16816 31340
rect 18788 31288 18840 31340
rect 13544 31220 13596 31272
rect 15476 31220 15528 31272
rect 17776 31220 17828 31272
rect 19708 31424 19760 31476
rect 25504 31424 25556 31476
rect 20168 31356 20220 31408
rect 21732 31356 21784 31408
rect 22008 31356 22060 31408
rect 22652 31356 22704 31408
rect 23020 31356 23072 31408
rect 20260 31288 20312 31340
rect 21456 31288 21508 31340
rect 13452 31127 13504 31136
rect 13452 31093 13461 31127
rect 13461 31093 13495 31127
rect 13495 31093 13504 31127
rect 13452 31084 13504 31093
rect 14464 31084 14516 31136
rect 16580 31084 16632 31136
rect 16856 31084 16908 31136
rect 17316 31084 17368 31136
rect 17684 31084 17736 31136
rect 18788 31084 18840 31136
rect 22468 31331 22520 31340
rect 22468 31297 22477 31331
rect 22477 31297 22511 31331
rect 22511 31297 22520 31331
rect 22468 31288 22520 31297
rect 24032 31288 24084 31340
rect 22376 31084 22428 31136
rect 23756 31084 23808 31136
rect 25504 31288 25556 31340
rect 24676 31084 24728 31136
rect 25136 31127 25188 31136
rect 25136 31093 25145 31127
rect 25145 31093 25179 31127
rect 25179 31093 25188 31127
rect 25136 31084 25188 31093
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 10232 30880 10284 30932
rect 8760 30676 8812 30728
rect 15292 30719 15344 30728
rect 15292 30685 15301 30719
rect 15301 30685 15335 30719
rect 15335 30685 15344 30719
rect 16304 30880 16356 30932
rect 17132 30880 17184 30932
rect 22652 30880 22704 30932
rect 25504 30923 25556 30932
rect 25504 30889 25513 30923
rect 25513 30889 25547 30923
rect 25547 30889 25556 30923
rect 25504 30880 25556 30889
rect 19432 30744 19484 30796
rect 22376 30744 22428 30796
rect 22652 30744 22704 30796
rect 15292 30676 15344 30685
rect 14832 30608 14884 30660
rect 20904 30608 20956 30660
rect 18328 30540 18380 30592
rect 18420 30540 18472 30592
rect 18788 30583 18840 30592
rect 18788 30549 18797 30583
rect 18797 30549 18831 30583
rect 18831 30549 18840 30583
rect 18788 30540 18840 30549
rect 20260 30583 20312 30592
rect 20260 30549 20269 30583
rect 20269 30549 20303 30583
rect 20303 30549 20312 30583
rect 20260 30540 20312 30549
rect 22376 30608 22428 30660
rect 24676 30540 24728 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 20260 30379 20312 30388
rect 20260 30345 20269 30379
rect 20269 30345 20303 30379
rect 20303 30345 20312 30379
rect 20260 30336 20312 30345
rect 11520 30268 11572 30320
rect 11888 30268 11940 30320
rect 15292 30268 15344 30320
rect 8576 30200 8628 30252
rect 13544 30243 13596 30252
rect 13544 30209 13553 30243
rect 13553 30209 13587 30243
rect 13587 30209 13596 30243
rect 13544 30200 13596 30209
rect 12808 30132 12860 30184
rect 13636 30132 13688 30184
rect 14556 30132 14608 30184
rect 19984 30268 20036 30320
rect 20536 30268 20588 30320
rect 16948 30200 17000 30252
rect 22192 30268 22244 30320
rect 22744 30268 22796 30320
rect 15568 30175 15620 30184
rect 15568 30141 15577 30175
rect 15577 30141 15611 30175
rect 15611 30141 15620 30175
rect 15568 30132 15620 30141
rect 16764 30175 16816 30184
rect 16764 30141 16773 30175
rect 16773 30141 16807 30175
rect 16807 30141 16816 30175
rect 24676 30200 24728 30252
rect 16764 30132 16816 30141
rect 20444 30175 20496 30184
rect 20444 30141 20453 30175
rect 20453 30141 20487 30175
rect 20487 30141 20496 30175
rect 20444 30132 20496 30141
rect 22560 30175 22612 30184
rect 22560 30141 22569 30175
rect 22569 30141 22603 30175
rect 22603 30141 22612 30175
rect 22560 30132 22612 30141
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 23664 30132 23716 30184
rect 24860 30132 24912 30184
rect 9036 30064 9088 30116
rect 16304 30064 16356 30116
rect 11796 30039 11848 30048
rect 11796 30005 11805 30039
rect 11805 30005 11839 30039
rect 11839 30005 11848 30039
rect 11796 29996 11848 30005
rect 15936 29996 15988 30048
rect 16948 30039 17000 30048
rect 16948 30005 16957 30039
rect 16957 30005 16991 30039
rect 16991 30005 17000 30039
rect 16948 29996 17000 30005
rect 18328 29996 18380 30048
rect 18788 29996 18840 30048
rect 20076 29996 20128 30048
rect 21732 29996 21784 30048
rect 26516 29996 26568 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 12808 29792 12860 29844
rect 12992 29792 13044 29844
rect 13452 29835 13504 29844
rect 13452 29801 13461 29835
rect 13461 29801 13495 29835
rect 13495 29801 13504 29835
rect 13452 29792 13504 29801
rect 16304 29835 16356 29844
rect 16304 29801 16313 29835
rect 16313 29801 16347 29835
rect 16347 29801 16356 29835
rect 16304 29792 16356 29801
rect 16948 29792 17000 29844
rect 22100 29792 22152 29844
rect 24584 29835 24636 29844
rect 24584 29801 24593 29835
rect 24593 29801 24627 29835
rect 24627 29801 24636 29835
rect 24584 29792 24636 29801
rect 11428 29656 11480 29708
rect 13636 29656 13688 29708
rect 15568 29724 15620 29776
rect 18972 29724 19024 29776
rect 23388 29724 23440 29776
rect 15844 29656 15896 29708
rect 19340 29656 19392 29708
rect 20352 29656 20404 29708
rect 15200 29588 15252 29640
rect 16304 29588 16356 29640
rect 20444 29588 20496 29640
rect 11060 29520 11112 29572
rect 11888 29520 11940 29572
rect 16580 29520 16632 29572
rect 18880 29520 18932 29572
rect 24492 29588 24544 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 24860 29520 24912 29572
rect 12716 29452 12768 29504
rect 16028 29452 16080 29504
rect 18420 29452 18472 29504
rect 19156 29452 19208 29504
rect 19984 29452 20036 29504
rect 22468 29452 22520 29504
rect 24032 29495 24084 29504
rect 24032 29461 24041 29495
rect 24041 29461 24075 29495
rect 24075 29461 24084 29495
rect 24032 29452 24084 29461
rect 24492 29495 24544 29504
rect 24492 29461 24501 29495
rect 24501 29461 24535 29495
rect 24535 29461 24544 29495
rect 24492 29452 24544 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 8852 29248 8904 29300
rect 12532 29291 12584 29300
rect 12532 29257 12541 29291
rect 12541 29257 12575 29291
rect 12575 29257 12584 29291
rect 12532 29248 12584 29257
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 13544 29248 13596 29300
rect 10232 29180 10284 29232
rect 10416 29112 10468 29164
rect 13636 29180 13688 29232
rect 15108 29291 15160 29300
rect 15108 29257 15117 29291
rect 15117 29257 15151 29291
rect 15151 29257 15160 29291
rect 15108 29248 15160 29257
rect 15936 29291 15988 29300
rect 15936 29257 15945 29291
rect 15945 29257 15979 29291
rect 15979 29257 15988 29291
rect 15936 29248 15988 29257
rect 16028 29291 16080 29300
rect 16028 29257 16037 29291
rect 16037 29257 16071 29291
rect 16071 29257 16080 29291
rect 16028 29248 16080 29257
rect 17408 29248 17460 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 19248 29291 19300 29300
rect 19248 29257 19257 29291
rect 19257 29257 19291 29291
rect 19291 29257 19300 29291
rect 19248 29248 19300 29257
rect 19340 29248 19392 29300
rect 23572 29248 23624 29300
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 9680 29044 9732 29096
rect 11520 29044 11572 29096
rect 12992 29044 13044 29096
rect 11980 28976 12032 29028
rect 11336 28908 11388 28960
rect 11796 28908 11848 28960
rect 14648 28976 14700 29028
rect 15752 28976 15804 29028
rect 19984 29223 20036 29232
rect 19984 29189 19993 29223
rect 19993 29189 20027 29223
rect 20027 29189 20036 29223
rect 19984 29180 20036 29189
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 19064 29044 19116 29096
rect 21272 29112 21324 29164
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 24584 29248 24636 29300
rect 25320 29248 25372 29300
rect 24952 29180 25004 29232
rect 25504 29180 25556 29232
rect 26424 29112 26476 29164
rect 23296 29044 23348 29096
rect 23480 29044 23532 29096
rect 23756 29044 23808 29096
rect 24952 29087 25004 29096
rect 24952 29053 24961 29087
rect 24961 29053 24995 29087
rect 24995 29053 25004 29087
rect 24952 29044 25004 29053
rect 17684 28976 17736 29028
rect 18788 29019 18840 29028
rect 18788 28985 18797 29019
rect 18797 28985 18831 29019
rect 18831 28985 18840 29019
rect 18788 28976 18840 28985
rect 24216 28976 24268 29028
rect 25872 28976 25924 29028
rect 26424 28976 26476 29028
rect 13360 28908 13412 28960
rect 16488 28908 16540 28960
rect 26884 28908 26936 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 9588 28704 9640 28756
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 23756 28704 23808 28756
rect 21916 28636 21968 28688
rect 22928 28636 22980 28688
rect 25872 28636 25924 28688
rect 15384 28611 15436 28620
rect 15384 28577 15393 28611
rect 15393 28577 15427 28611
rect 15427 28577 15436 28611
rect 15384 28568 15436 28577
rect 15476 28568 15528 28620
rect 16396 28568 16448 28620
rect 18696 28568 18748 28620
rect 20904 28568 20956 28620
rect 21364 28568 21416 28620
rect 11428 28543 11480 28552
rect 11428 28509 11437 28543
rect 11437 28509 11471 28543
rect 11471 28509 11480 28543
rect 11428 28500 11480 28509
rect 14832 28500 14884 28552
rect 20444 28500 20496 28552
rect 22100 28568 22152 28620
rect 25412 28568 25464 28620
rect 23940 28500 23992 28552
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 25228 28500 25280 28552
rect 9588 28432 9640 28484
rect 10968 28432 11020 28484
rect 11336 28432 11388 28484
rect 12716 28432 12768 28484
rect 16396 28432 16448 28484
rect 13360 28364 13412 28416
rect 13544 28407 13596 28416
rect 13544 28373 13553 28407
rect 13553 28373 13587 28407
rect 13587 28373 13596 28407
rect 13544 28364 13596 28373
rect 13820 28364 13872 28416
rect 15568 28364 15620 28416
rect 16120 28407 16172 28416
rect 16120 28373 16129 28407
rect 16129 28373 16163 28407
rect 16163 28373 16172 28407
rect 16120 28364 16172 28373
rect 16304 28407 16356 28416
rect 16304 28373 16313 28407
rect 16313 28373 16347 28407
rect 16347 28373 16356 28407
rect 16304 28364 16356 28373
rect 19064 28432 19116 28484
rect 21364 28432 21416 28484
rect 26056 28432 26108 28484
rect 18328 28364 18380 28416
rect 19524 28364 19576 28416
rect 19800 28407 19852 28416
rect 19800 28373 19809 28407
rect 19809 28373 19843 28407
rect 19843 28373 19852 28407
rect 19800 28364 19852 28373
rect 21640 28364 21692 28416
rect 22192 28364 22244 28416
rect 22652 28364 22704 28416
rect 23940 28407 23992 28416
rect 23940 28373 23949 28407
rect 23949 28373 23983 28407
rect 23983 28373 23992 28407
rect 23940 28364 23992 28373
rect 24400 28364 24452 28416
rect 24492 28364 24544 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 12716 28160 12768 28212
rect 13544 28160 13596 28212
rect 16396 28160 16448 28212
rect 16672 28092 16724 28144
rect 18604 28092 18656 28144
rect 19800 28160 19852 28212
rect 26240 28160 26292 28212
rect 16488 28024 16540 28076
rect 17316 28067 17368 28076
rect 17316 28033 17325 28067
rect 17325 28033 17359 28067
rect 17359 28033 17368 28067
rect 17316 28024 17368 28033
rect 18512 28024 18564 28076
rect 9864 27888 9916 27940
rect 12072 27956 12124 28008
rect 13452 27956 13504 28008
rect 15384 27956 15436 28008
rect 14832 27888 14884 27940
rect 17408 27999 17460 28008
rect 17408 27965 17417 27999
rect 17417 27965 17451 27999
rect 17451 27965 17460 27999
rect 17408 27956 17460 27965
rect 17960 27956 18012 28008
rect 18328 27956 18380 28008
rect 20444 27999 20496 28008
rect 20444 27965 20453 27999
rect 20453 27965 20487 27999
rect 20487 27965 20496 27999
rect 20444 27956 20496 27965
rect 20812 28092 20864 28144
rect 21364 28092 21416 28144
rect 21548 28092 21600 28144
rect 22560 28092 22612 28144
rect 22928 28092 22980 28144
rect 24400 28092 24452 28144
rect 24676 28092 24728 28144
rect 24952 28092 25004 28144
rect 21272 28067 21324 28076
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 16672 27888 16724 27940
rect 17040 27888 17092 27940
rect 21272 27888 21324 27940
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 24124 27956 24176 28008
rect 24676 27999 24728 28008
rect 24676 27965 24685 27999
rect 24685 27965 24719 27999
rect 24719 27965 24728 27999
rect 24676 27956 24728 27965
rect 13452 27863 13504 27872
rect 13452 27829 13461 27863
rect 13461 27829 13495 27863
rect 13495 27829 13504 27863
rect 13452 27820 13504 27829
rect 13912 27820 13964 27872
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 18512 27863 18564 27872
rect 18512 27829 18521 27863
rect 18521 27829 18555 27863
rect 18555 27829 18564 27863
rect 18512 27820 18564 27829
rect 18604 27820 18656 27872
rect 21548 27863 21600 27872
rect 21548 27829 21557 27863
rect 21557 27829 21591 27863
rect 21591 27829 21600 27863
rect 21548 27820 21600 27829
rect 21640 27820 21692 27872
rect 22744 27820 22796 27872
rect 23388 27820 23440 27872
rect 23572 27820 23624 27872
rect 25412 27863 25464 27872
rect 25412 27829 25421 27863
rect 25421 27829 25455 27863
rect 25455 27829 25464 27863
rect 25412 27820 25464 27829
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 13452 27616 13504 27668
rect 22100 27659 22152 27668
rect 22100 27625 22109 27659
rect 22109 27625 22143 27659
rect 22143 27625 22152 27659
rect 22100 27616 22152 27625
rect 23388 27616 23440 27668
rect 12348 27548 12400 27600
rect 12716 27548 12768 27600
rect 24676 27548 24728 27600
rect 11428 27480 11480 27532
rect 11244 27344 11296 27396
rect 9312 27276 9364 27328
rect 16212 27480 16264 27532
rect 17776 27480 17828 27532
rect 23572 27480 23624 27532
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 12716 27412 12768 27464
rect 13820 27412 13872 27464
rect 14924 27412 14976 27464
rect 16764 27412 16816 27464
rect 17960 27412 18012 27464
rect 13912 27344 13964 27396
rect 20812 27344 20864 27396
rect 22008 27344 22060 27396
rect 24860 27412 24912 27464
rect 25412 27412 25464 27464
rect 12624 27276 12676 27328
rect 13544 27276 13596 27328
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 16120 27276 16172 27328
rect 16304 27276 16356 27328
rect 16488 27276 16540 27328
rect 17592 27276 17644 27328
rect 20720 27276 20772 27328
rect 22652 27276 22704 27328
rect 26056 27344 26108 27396
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 9588 27072 9640 27124
rect 9864 27004 9916 27056
rect 11060 27115 11112 27124
rect 11060 27081 11069 27115
rect 11069 27081 11103 27115
rect 11103 27081 11112 27115
rect 11060 27072 11112 27081
rect 16856 27072 16908 27124
rect 11244 27004 11296 27056
rect 12716 27004 12768 27056
rect 15108 27004 15160 27056
rect 15752 27047 15804 27056
rect 15752 27013 15761 27047
rect 15761 27013 15795 27047
rect 15795 27013 15804 27047
rect 15752 27004 15804 27013
rect 15936 27004 15988 27056
rect 21548 27072 21600 27124
rect 22376 27072 22428 27124
rect 22836 27115 22888 27124
rect 22836 27081 22845 27115
rect 22845 27081 22879 27115
rect 22879 27081 22888 27115
rect 22836 27072 22888 27081
rect 22100 27004 22152 27056
rect 22560 27004 22612 27056
rect 14832 26979 14884 26988
rect 14832 26945 14841 26979
rect 14841 26945 14875 26979
rect 14875 26945 14884 26979
rect 14832 26936 14884 26945
rect 18328 26936 18380 26988
rect 22192 26936 22244 26988
rect 22376 26936 22428 26988
rect 9312 26800 9364 26852
rect 11244 26732 11296 26784
rect 12348 26732 12400 26784
rect 12532 26732 12584 26784
rect 15016 26732 15068 26784
rect 18696 26732 18748 26784
rect 19432 26732 19484 26784
rect 20444 26868 20496 26920
rect 23664 27072 23716 27124
rect 24676 27072 24728 27124
rect 24952 26936 25004 26988
rect 23572 26911 23624 26920
rect 23572 26877 23581 26911
rect 23581 26877 23615 26911
rect 23615 26877 23624 26911
rect 23572 26868 23624 26877
rect 25412 26868 25464 26920
rect 21272 26800 21324 26852
rect 20168 26732 20220 26784
rect 20812 26732 20864 26784
rect 22008 26775 22060 26784
rect 22008 26741 22017 26775
rect 22017 26741 22051 26775
rect 22051 26741 22060 26775
rect 22008 26732 22060 26741
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 9404 26528 9456 26580
rect 12072 26528 12124 26580
rect 13636 26528 13688 26580
rect 16396 26528 16448 26580
rect 17224 26571 17276 26580
rect 17224 26537 17233 26571
rect 17233 26537 17267 26571
rect 17267 26537 17276 26571
rect 17224 26528 17276 26537
rect 22100 26528 22152 26580
rect 24952 26528 25004 26580
rect 11520 26460 11572 26512
rect 11612 26460 11664 26512
rect 9864 26392 9916 26444
rect 14740 26392 14792 26444
rect 15476 26392 15528 26444
rect 16580 26460 16632 26512
rect 17132 26460 17184 26512
rect 20812 26460 20864 26512
rect 22560 26460 22612 26512
rect 25228 26460 25280 26512
rect 16212 26435 16264 26444
rect 16212 26401 16221 26435
rect 16221 26401 16255 26435
rect 16255 26401 16264 26435
rect 16212 26392 16264 26401
rect 16764 26435 16816 26444
rect 16764 26401 16773 26435
rect 16773 26401 16807 26435
rect 16807 26401 16816 26435
rect 16764 26392 16816 26401
rect 16948 26435 17000 26444
rect 16948 26401 16957 26435
rect 16957 26401 16991 26435
rect 16991 26401 17000 26435
rect 16948 26392 17000 26401
rect 20720 26392 20772 26444
rect 22284 26392 22336 26444
rect 25044 26392 25096 26444
rect 13452 26324 13504 26376
rect 8484 26256 8536 26308
rect 9404 26299 9456 26308
rect 9404 26265 9413 26299
rect 9413 26265 9447 26299
rect 9447 26265 9456 26299
rect 9404 26256 9456 26265
rect 11244 26299 11296 26308
rect 11244 26265 11253 26299
rect 11253 26265 11287 26299
rect 11287 26265 11296 26299
rect 11244 26256 11296 26265
rect 14924 26188 14976 26240
rect 16396 26256 16448 26308
rect 18328 26324 18380 26376
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 23296 26324 23348 26376
rect 23848 26367 23900 26376
rect 23848 26333 23857 26367
rect 23857 26333 23891 26367
rect 23891 26333 23900 26367
rect 23848 26324 23900 26333
rect 17316 26256 17368 26308
rect 20168 26256 20220 26308
rect 22376 26299 22428 26308
rect 22376 26265 22385 26299
rect 22385 26265 22419 26299
rect 22419 26265 22428 26299
rect 22376 26256 22428 26265
rect 26056 26324 26108 26376
rect 25136 26256 25188 26308
rect 18328 26188 18380 26240
rect 25872 26188 25924 26240
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 12624 25984 12676 26036
rect 16856 25984 16908 26036
rect 18328 25984 18380 26036
rect 19064 25984 19116 26036
rect 22192 25984 22244 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 11428 25916 11480 25968
rect 9956 25848 10008 25900
rect 14648 25848 14700 25900
rect 18972 25916 19024 25968
rect 11060 25780 11112 25832
rect 13360 25780 13412 25832
rect 15384 25823 15436 25832
rect 15384 25789 15393 25823
rect 15393 25789 15427 25823
rect 15427 25789 15436 25823
rect 15384 25780 15436 25789
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 21456 25848 21508 25900
rect 24768 25984 24820 26036
rect 24860 25916 24912 25968
rect 23940 25891 23992 25900
rect 23940 25857 23949 25891
rect 23949 25857 23983 25891
rect 23983 25857 23992 25891
rect 23940 25848 23992 25857
rect 17408 25823 17460 25832
rect 17408 25789 17417 25823
rect 17417 25789 17451 25823
rect 17451 25789 17460 25823
rect 17408 25780 17460 25789
rect 13820 25644 13872 25696
rect 17592 25712 17644 25764
rect 18420 25823 18472 25832
rect 18420 25789 18429 25823
rect 18429 25789 18463 25823
rect 18463 25789 18472 25823
rect 18420 25780 18472 25789
rect 20904 25780 20956 25832
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 17040 25687 17092 25696
rect 17040 25653 17049 25687
rect 17049 25653 17083 25687
rect 17083 25653 17092 25687
rect 17040 25644 17092 25653
rect 17408 25644 17460 25696
rect 18328 25644 18380 25696
rect 19064 25687 19116 25696
rect 19064 25653 19073 25687
rect 19073 25653 19107 25687
rect 19107 25653 19116 25687
rect 19064 25644 19116 25653
rect 21456 25644 21508 25696
rect 22008 25687 22060 25696
rect 22008 25653 22017 25687
rect 22017 25653 22051 25687
rect 22051 25653 22060 25687
rect 22008 25644 22060 25653
rect 25596 25712 25648 25764
rect 23388 25644 23440 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 11704 25440 11756 25492
rect 21548 25440 21600 25492
rect 23940 25440 23992 25492
rect 24860 25440 24912 25492
rect 25596 25440 25648 25492
rect 25780 25440 25832 25492
rect 14648 25372 14700 25424
rect 15200 25372 15252 25424
rect 14740 25304 14792 25356
rect 11244 25236 11296 25288
rect 12808 25236 12860 25288
rect 9680 25100 9732 25152
rect 10784 25100 10836 25152
rect 14832 25168 14884 25220
rect 12900 25100 12952 25152
rect 12992 25143 13044 25152
rect 12992 25109 13001 25143
rect 13001 25109 13035 25143
rect 13035 25109 13044 25143
rect 12992 25100 13044 25109
rect 14648 25143 14700 25152
rect 14648 25109 14657 25143
rect 14657 25109 14691 25143
rect 14691 25109 14700 25143
rect 14648 25100 14700 25109
rect 15844 25168 15896 25220
rect 18604 25372 18656 25424
rect 19892 25372 19944 25424
rect 20352 25415 20404 25424
rect 20352 25381 20361 25415
rect 20361 25381 20395 25415
rect 20395 25381 20404 25415
rect 20352 25372 20404 25381
rect 17040 25304 17092 25356
rect 16948 25279 17000 25288
rect 16948 25245 16957 25279
rect 16957 25245 16991 25279
rect 16991 25245 17000 25279
rect 16948 25236 17000 25245
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 15292 25143 15344 25152
rect 15292 25109 15301 25143
rect 15301 25109 15335 25143
rect 15335 25109 15344 25143
rect 15292 25100 15344 25109
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 16304 25100 16356 25152
rect 18328 25236 18380 25288
rect 20352 25236 20404 25288
rect 18328 25143 18380 25152
rect 18328 25109 18337 25143
rect 18337 25109 18371 25143
rect 18371 25109 18380 25143
rect 18328 25100 18380 25109
rect 18512 25100 18564 25152
rect 19708 25211 19760 25220
rect 19708 25177 19717 25211
rect 19717 25177 19751 25211
rect 19751 25177 19760 25211
rect 19708 25168 19760 25177
rect 23848 25372 23900 25424
rect 24676 25372 24728 25424
rect 21548 25279 21600 25288
rect 21548 25245 21557 25279
rect 21557 25245 21591 25279
rect 21591 25245 21600 25279
rect 21548 25236 21600 25245
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 23848 25211 23900 25220
rect 23848 25177 23857 25211
rect 23857 25177 23891 25211
rect 23891 25177 23900 25211
rect 23848 25168 23900 25177
rect 22192 25100 22244 25152
rect 25504 25100 25556 25152
rect 25872 25100 25924 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 10508 24896 10560 24948
rect 15292 24896 15344 24948
rect 17224 24939 17276 24948
rect 17224 24905 17233 24939
rect 17233 24905 17267 24939
rect 17267 24905 17276 24939
rect 17224 24896 17276 24905
rect 19892 24896 19944 24948
rect 11796 24828 11848 24880
rect 12716 24828 12768 24880
rect 12992 24828 13044 24880
rect 18604 24828 18656 24880
rect 9128 24760 9180 24812
rect 11980 24803 12032 24812
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 11980 24760 12032 24769
rect 14832 24760 14884 24812
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 15844 24760 15896 24812
rect 11152 24735 11204 24744
rect 11152 24701 11161 24735
rect 11161 24701 11195 24735
rect 11195 24701 11204 24735
rect 11152 24692 11204 24701
rect 12072 24692 12124 24744
rect 12900 24692 12952 24744
rect 13452 24692 13504 24744
rect 13728 24692 13780 24744
rect 9404 24599 9456 24608
rect 9404 24565 9413 24599
rect 9413 24565 9447 24599
rect 9447 24565 9456 24599
rect 9404 24556 9456 24565
rect 11060 24556 11112 24608
rect 16948 24692 17000 24744
rect 17040 24692 17092 24744
rect 18328 24760 18380 24812
rect 20260 24828 20312 24880
rect 24124 24828 24176 24880
rect 18420 24692 18472 24744
rect 15384 24624 15436 24676
rect 22652 24760 22704 24812
rect 24952 24760 25004 24812
rect 19156 24692 19208 24744
rect 19432 24692 19484 24744
rect 20076 24692 20128 24744
rect 22284 24692 22336 24744
rect 22744 24735 22796 24744
rect 22744 24701 22753 24735
rect 22753 24701 22787 24735
rect 22787 24701 22796 24735
rect 22744 24692 22796 24701
rect 23296 24692 23348 24744
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 25044 24692 25096 24744
rect 25412 24692 25464 24744
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 16488 24556 16540 24608
rect 21548 24624 21600 24676
rect 18328 24556 18380 24608
rect 18420 24556 18472 24608
rect 19708 24556 19760 24608
rect 21364 24556 21416 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 9404 24352 9456 24404
rect 9588 24352 9640 24404
rect 13728 24395 13780 24404
rect 13728 24361 13737 24395
rect 13737 24361 13771 24395
rect 13771 24361 13780 24395
rect 13728 24352 13780 24361
rect 14740 24284 14792 24336
rect 18880 24284 18932 24336
rect 11152 24216 11204 24268
rect 12348 24216 12400 24268
rect 12716 24216 12768 24268
rect 15476 24216 15528 24268
rect 18696 24259 18748 24268
rect 18696 24225 18705 24259
rect 18705 24225 18739 24259
rect 18739 24225 18748 24259
rect 18696 24216 18748 24225
rect 7840 24148 7892 24200
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 21640 24352 21692 24404
rect 24952 24352 25004 24404
rect 25136 24352 25188 24404
rect 25320 24352 25372 24404
rect 23296 24284 23348 24336
rect 19156 24216 19208 24268
rect 24124 24216 24176 24268
rect 9496 24080 9548 24132
rect 11244 24123 11296 24132
rect 8392 24012 8444 24064
rect 9128 24012 9180 24064
rect 11244 24089 11253 24123
rect 11253 24089 11287 24123
rect 11287 24089 11296 24123
rect 11244 24080 11296 24089
rect 11520 24080 11572 24132
rect 12532 24080 12584 24132
rect 12716 24080 12768 24132
rect 18972 24080 19024 24132
rect 20352 24080 20404 24132
rect 20444 24080 20496 24132
rect 11152 24012 11204 24064
rect 16672 24012 16724 24064
rect 16764 24012 16816 24064
rect 18512 24012 18564 24064
rect 20076 24012 20128 24064
rect 20904 24123 20956 24132
rect 20904 24089 20913 24123
rect 20913 24089 20947 24123
rect 20947 24089 20956 24123
rect 20904 24080 20956 24089
rect 22284 24080 22336 24132
rect 21548 24055 21600 24064
rect 21548 24021 21557 24055
rect 21557 24021 21591 24055
rect 21591 24021 21600 24055
rect 21548 24012 21600 24021
rect 23480 24012 23532 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 8392 23740 8444 23792
rect 10416 23851 10468 23860
rect 10416 23817 10425 23851
rect 10425 23817 10459 23851
rect 10459 23817 10468 23851
rect 10416 23808 10468 23817
rect 13360 23808 13412 23860
rect 13636 23783 13688 23792
rect 13636 23749 13645 23783
rect 13645 23749 13679 23783
rect 13679 23749 13688 23783
rect 13636 23740 13688 23749
rect 13728 23740 13780 23792
rect 15016 23808 15068 23860
rect 16764 23808 16816 23860
rect 17500 23808 17552 23860
rect 17868 23808 17920 23860
rect 14924 23740 14976 23792
rect 13544 23672 13596 23724
rect 7840 23604 7892 23656
rect 10508 23604 10560 23656
rect 10876 23647 10928 23656
rect 10876 23613 10885 23647
rect 10885 23613 10919 23647
rect 10919 23613 10928 23647
rect 10876 23604 10928 23613
rect 10968 23647 11020 23656
rect 10968 23613 10977 23647
rect 10977 23613 11011 23647
rect 11011 23613 11020 23647
rect 10968 23604 11020 23613
rect 13452 23604 13504 23656
rect 10784 23468 10836 23520
rect 12532 23468 12584 23520
rect 13544 23468 13596 23520
rect 17040 23672 17092 23724
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 18512 23783 18564 23792
rect 18512 23749 18521 23783
rect 18521 23749 18555 23783
rect 18555 23749 18564 23783
rect 18512 23740 18564 23749
rect 19248 23740 19300 23792
rect 21916 23808 21968 23860
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 20260 23740 20312 23792
rect 20720 23740 20772 23792
rect 19984 23604 20036 23656
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 20904 23604 20956 23656
rect 21548 23783 21600 23792
rect 21548 23749 21557 23783
rect 21557 23749 21591 23783
rect 21591 23749 21600 23783
rect 25044 23808 25096 23860
rect 21548 23740 21600 23749
rect 25136 23740 25188 23792
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 23204 23647 23256 23656
rect 23204 23613 23213 23647
rect 23213 23613 23247 23647
rect 23247 23613 23256 23647
rect 23204 23604 23256 23613
rect 23480 23647 23532 23656
rect 23480 23613 23489 23647
rect 23489 23613 23523 23647
rect 23523 23613 23532 23647
rect 23480 23604 23532 23613
rect 17132 23468 17184 23520
rect 17316 23468 17368 23520
rect 17500 23468 17552 23520
rect 18144 23468 18196 23520
rect 18420 23468 18472 23520
rect 18972 23511 19024 23520
rect 18972 23477 18981 23511
rect 18981 23477 19015 23511
rect 19015 23477 19024 23511
rect 18972 23468 19024 23477
rect 19800 23536 19852 23588
rect 21916 23468 21968 23520
rect 23940 23468 23992 23520
rect 25136 23468 25188 23520
rect 25504 23468 25556 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 9220 23264 9272 23316
rect 10508 23264 10560 23316
rect 11060 23264 11112 23316
rect 11336 23264 11388 23316
rect 11888 23264 11940 23316
rect 8208 23196 8260 23248
rect 8668 23128 8720 23180
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 12992 23128 13044 23180
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 10416 22992 10468 23044
rect 11336 22992 11388 23044
rect 15660 23060 15712 23112
rect 10048 22924 10100 22976
rect 11244 22967 11296 22976
rect 11244 22933 11253 22967
rect 11253 22933 11287 22967
rect 11287 22933 11296 22967
rect 11244 22924 11296 22933
rect 12624 22924 12676 22976
rect 14464 22924 14516 22976
rect 17316 23264 17368 23316
rect 19432 23196 19484 23248
rect 25504 23264 25556 23316
rect 26056 23264 26108 23316
rect 26424 23196 26476 23248
rect 18420 23128 18472 23180
rect 19064 23128 19116 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 20812 23128 20864 23180
rect 24860 23128 24912 23180
rect 24952 23128 25004 23180
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 18604 23060 18656 23112
rect 20260 23060 20312 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 24032 23060 24084 23112
rect 17868 22924 17920 22976
rect 18512 22992 18564 23044
rect 18696 22924 18748 22976
rect 22008 22992 22060 23044
rect 25136 22992 25188 23044
rect 22100 22924 22152 22976
rect 24032 22924 24084 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 7564 22720 7616 22772
rect 8300 22720 8352 22772
rect 9588 22695 9640 22704
rect 9588 22661 9597 22695
rect 9597 22661 9631 22695
rect 9631 22661 9640 22695
rect 9588 22652 9640 22661
rect 9680 22652 9732 22704
rect 12808 22720 12860 22772
rect 8300 22584 8352 22636
rect 12716 22652 12768 22704
rect 14464 22763 14516 22772
rect 14464 22729 14473 22763
rect 14473 22729 14507 22763
rect 14507 22729 14516 22763
rect 14464 22720 14516 22729
rect 14832 22720 14884 22772
rect 18604 22720 18656 22772
rect 19616 22720 19668 22772
rect 24676 22720 24728 22772
rect 21640 22652 21692 22704
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 13912 22584 13964 22636
rect 18696 22584 18748 22636
rect 20444 22584 20496 22636
rect 21456 22584 21508 22636
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 23940 22627 23992 22636
rect 23940 22593 23949 22627
rect 23949 22593 23983 22627
rect 23983 22593 23992 22627
rect 23940 22584 23992 22593
rect 19708 22516 19760 22568
rect 22836 22559 22888 22568
rect 22836 22525 22845 22559
rect 22845 22525 22879 22559
rect 22879 22525 22888 22559
rect 22836 22516 22888 22525
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 9404 22380 9456 22432
rect 18604 22448 18656 22500
rect 20812 22448 20864 22500
rect 12992 22380 13044 22432
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 9772 22176 9824 22228
rect 15936 22176 15988 22228
rect 18696 22176 18748 22228
rect 21088 22176 21140 22228
rect 23848 22176 23900 22228
rect 6920 22108 6972 22160
rect 7840 22108 7892 22160
rect 9680 22108 9732 22160
rect 11060 22108 11112 22160
rect 11152 22108 11204 22160
rect 12532 22108 12584 22160
rect 14096 22040 14148 22092
rect 14556 22040 14608 22092
rect 15752 22108 15804 22160
rect 17868 22108 17920 22160
rect 16948 22040 17000 22092
rect 19064 22040 19116 22092
rect 20628 22040 20680 22092
rect 25412 22176 25464 22228
rect 21548 21972 21600 22024
rect 23296 22015 23348 22024
rect 23296 21981 23305 22015
rect 23305 21981 23339 22015
rect 23339 21981 23348 22015
rect 23296 21972 23348 21981
rect 11152 21904 11204 21956
rect 15936 21904 15988 21956
rect 16488 21904 16540 21956
rect 8300 21836 8352 21888
rect 10600 21836 10652 21888
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 11428 21879 11480 21888
rect 11428 21845 11437 21879
rect 11437 21845 11471 21879
rect 11471 21845 11480 21879
rect 11428 21836 11480 21845
rect 13912 21836 13964 21888
rect 14004 21836 14056 21888
rect 15844 21836 15896 21888
rect 17408 21836 17460 21888
rect 23020 21947 23072 21956
rect 23020 21913 23029 21947
rect 23029 21913 23063 21947
rect 23063 21913 23072 21947
rect 23020 21904 23072 21913
rect 17868 21879 17920 21888
rect 17868 21845 17877 21879
rect 17877 21845 17911 21879
rect 17911 21845 17920 21879
rect 17868 21836 17920 21845
rect 19616 21836 19668 21888
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 20352 21836 20404 21888
rect 20904 21836 20956 21888
rect 22008 21836 22060 21888
rect 25228 21972 25280 22024
rect 24400 21836 24452 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 8668 21675 8720 21684
rect 8668 21641 8677 21675
rect 8677 21641 8711 21675
rect 8711 21641 8720 21675
rect 8668 21632 8720 21641
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 10232 21632 10284 21684
rect 11060 21632 11112 21684
rect 12716 21632 12768 21684
rect 12164 21564 12216 21616
rect 15108 21632 15160 21684
rect 18696 21632 18748 21684
rect 20076 21632 20128 21684
rect 22560 21632 22612 21684
rect 23296 21632 23348 21684
rect 14280 21564 14332 21616
rect 8300 21496 8352 21548
rect 9220 21496 9272 21548
rect 9956 21496 10008 21548
rect 11612 21496 11664 21548
rect 18788 21564 18840 21616
rect 19984 21564 20036 21616
rect 21548 21564 21600 21616
rect 15844 21496 15896 21548
rect 22192 21496 22244 21548
rect 6920 21471 6972 21480
rect 6920 21437 6929 21471
rect 6929 21437 6963 21471
rect 6963 21437 6972 21471
rect 6920 21428 6972 21437
rect 7748 21428 7800 21480
rect 9312 21471 9364 21480
rect 9312 21437 9321 21471
rect 9321 21437 9355 21471
rect 9355 21437 9364 21471
rect 9312 21428 9364 21437
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 19708 21471 19760 21480
rect 19708 21437 19717 21471
rect 19717 21437 19751 21471
rect 19751 21437 19760 21471
rect 19708 21428 19760 21437
rect 23480 21428 23532 21480
rect 23572 21428 23624 21480
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 21640 21360 21692 21412
rect 22836 21360 22888 21412
rect 24400 21428 24452 21480
rect 25320 21428 25372 21480
rect 12716 21292 12768 21344
rect 13544 21292 13596 21344
rect 15108 21335 15160 21344
rect 15108 21301 15117 21335
rect 15117 21301 15151 21335
rect 15151 21301 15160 21335
rect 15108 21292 15160 21301
rect 18788 21292 18840 21344
rect 20444 21292 20496 21344
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 23020 21292 23072 21344
rect 23296 21335 23348 21344
rect 23296 21301 23305 21335
rect 23305 21301 23339 21335
rect 23339 21301 23348 21335
rect 23296 21292 23348 21301
rect 24952 21292 25004 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 21088 21088 21140 21140
rect 9680 20952 9732 21004
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 12072 20884 12124 20936
rect 10968 20859 11020 20868
rect 10968 20825 10977 20859
rect 10977 20825 11011 20859
rect 11011 20825 11020 20859
rect 10968 20816 11020 20825
rect 12808 20816 12860 20868
rect 9220 20748 9272 20800
rect 12532 20748 12584 20800
rect 15200 20952 15252 21004
rect 16948 20995 17000 21004
rect 16948 20961 16957 20995
rect 16957 20961 16991 20995
rect 16991 20961 17000 20995
rect 16948 20952 17000 20961
rect 19616 20995 19668 21004
rect 19616 20961 19625 20995
rect 19625 20961 19659 20995
rect 19659 20961 19668 20995
rect 19616 20952 19668 20961
rect 17224 20884 17276 20936
rect 17776 20884 17828 20936
rect 19248 20884 19300 20936
rect 22192 20995 22244 21004
rect 22192 20961 22201 20995
rect 22201 20961 22235 20995
rect 22235 20961 22244 20995
rect 22192 20952 22244 20961
rect 24676 20995 24728 21004
rect 24676 20961 24685 20995
rect 24685 20961 24719 20995
rect 24719 20961 24728 20995
rect 24676 20952 24728 20961
rect 24952 20952 25004 21004
rect 25412 20952 25464 21004
rect 24860 20884 24912 20936
rect 25044 20884 25096 20936
rect 16580 20816 16632 20868
rect 19064 20816 19116 20868
rect 14648 20791 14700 20800
rect 14648 20757 14657 20791
rect 14657 20757 14691 20791
rect 14691 20757 14700 20791
rect 14648 20748 14700 20757
rect 15844 20748 15896 20800
rect 17224 20791 17276 20800
rect 17224 20757 17233 20791
rect 17233 20757 17267 20791
rect 17267 20757 17276 20791
rect 17224 20748 17276 20757
rect 17408 20748 17460 20800
rect 19892 20748 19944 20800
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 25044 20748 25096 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 8300 20476 8352 20528
rect 10416 20587 10468 20596
rect 10416 20553 10425 20587
rect 10425 20553 10459 20587
rect 10459 20553 10468 20587
rect 10416 20544 10468 20553
rect 11336 20544 11388 20596
rect 15384 20544 15436 20596
rect 16764 20544 16816 20596
rect 18420 20544 18472 20596
rect 14648 20476 14700 20528
rect 15108 20476 15160 20528
rect 6552 20408 6604 20460
rect 6920 20408 6972 20460
rect 12440 20408 12492 20460
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 17224 20408 17276 20460
rect 19156 20408 19208 20460
rect 20168 20476 20220 20528
rect 21732 20544 21784 20596
rect 23572 20544 23624 20596
rect 23848 20544 23900 20596
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 20812 20519 20864 20528
rect 20812 20485 20821 20519
rect 20821 20485 20855 20519
rect 20855 20485 20864 20519
rect 20812 20476 20864 20485
rect 21640 20476 21692 20528
rect 8668 20340 8720 20392
rect 10140 20340 10192 20392
rect 10416 20340 10468 20392
rect 10784 20272 10836 20324
rect 12716 20272 12768 20324
rect 17868 20340 17920 20392
rect 20536 20383 20588 20392
rect 20536 20349 20545 20383
rect 20545 20349 20579 20383
rect 20579 20349 20588 20383
rect 20536 20340 20588 20349
rect 21088 20340 21140 20392
rect 23572 20383 23624 20392
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 23572 20340 23624 20349
rect 25136 20340 25188 20392
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 16764 20204 16816 20256
rect 17040 20204 17092 20256
rect 23480 20272 23532 20324
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19708 20247 19760 20256
rect 19708 20213 19717 20247
rect 19717 20213 19751 20247
rect 19751 20213 19760 20247
rect 19708 20204 19760 20213
rect 21732 20204 21784 20256
rect 22744 20204 22796 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 10968 20000 11020 20052
rect 13360 20000 13412 20052
rect 15108 20000 15160 20052
rect 16580 20000 16632 20052
rect 17040 20000 17092 20052
rect 21180 20000 21232 20052
rect 23664 20000 23716 20052
rect 24676 20000 24728 20052
rect 17224 19932 17276 19984
rect 9404 19907 9456 19916
rect 9404 19873 9413 19907
rect 9413 19873 9447 19907
rect 9447 19873 9456 19907
rect 9404 19864 9456 19873
rect 11520 19907 11572 19916
rect 11520 19873 11529 19907
rect 11529 19873 11563 19907
rect 11563 19873 11572 19907
rect 11520 19864 11572 19873
rect 12440 19864 12492 19916
rect 13360 19864 13412 19916
rect 14280 19907 14332 19916
rect 14280 19873 14289 19907
rect 14289 19873 14323 19907
rect 14323 19873 14332 19907
rect 14280 19864 14332 19873
rect 14556 19864 14608 19916
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 17868 19864 17920 19916
rect 20260 19864 20312 19916
rect 18328 19796 18380 19848
rect 19524 19796 19576 19848
rect 8300 19660 8352 19712
rect 14832 19728 14884 19780
rect 15108 19728 15160 19780
rect 9588 19660 9640 19712
rect 11428 19660 11480 19712
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 16488 19660 16540 19712
rect 19800 19728 19852 19780
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 21548 19728 21600 19780
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 21640 19703 21692 19712
rect 21640 19669 21649 19703
rect 21649 19669 21683 19703
rect 21683 19669 21692 19703
rect 23848 19728 23900 19780
rect 24124 19771 24176 19780
rect 24124 19737 24133 19771
rect 24133 19737 24167 19771
rect 24167 19737 24176 19771
rect 24124 19728 24176 19737
rect 21640 19660 21692 19669
rect 24952 19660 25004 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 9588 19456 9640 19508
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 12440 19456 12492 19508
rect 15200 19499 15252 19508
rect 15200 19465 15209 19499
rect 15209 19465 15243 19499
rect 15243 19465 15252 19499
rect 15200 19456 15252 19465
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 19248 19456 19300 19508
rect 20444 19499 20496 19508
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 20720 19456 20772 19508
rect 22468 19456 22520 19508
rect 24032 19456 24084 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 8208 19388 8260 19440
rect 13912 19388 13964 19440
rect 14464 19388 14516 19440
rect 15752 19388 15804 19440
rect 9036 19320 9088 19372
rect 9956 19320 10008 19372
rect 14280 19363 14332 19372
rect 14280 19329 14289 19363
rect 14289 19329 14323 19363
rect 14323 19329 14332 19363
rect 14280 19320 14332 19329
rect 15016 19363 15068 19372
rect 15016 19329 15025 19363
rect 15025 19329 15059 19363
rect 15059 19329 15068 19363
rect 15016 19320 15068 19329
rect 16396 19320 16448 19372
rect 17040 19320 17092 19372
rect 20536 19320 20588 19372
rect 22100 19388 22152 19440
rect 23572 19388 23624 19440
rect 23664 19431 23716 19440
rect 23664 19397 23673 19431
rect 23673 19397 23707 19431
rect 23707 19397 23716 19431
rect 23664 19388 23716 19397
rect 24124 19388 24176 19440
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 6920 19252 6972 19304
rect 7564 19252 7616 19304
rect 8668 19252 8720 19304
rect 9404 19252 9456 19304
rect 7840 19184 7892 19236
rect 10784 19184 10836 19236
rect 11428 19184 11480 19236
rect 14648 19184 14700 19236
rect 16580 19252 16632 19304
rect 21640 19252 21692 19304
rect 23296 19252 23348 19304
rect 18788 19184 18840 19236
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 9588 19116 9640 19168
rect 13912 19116 13964 19168
rect 14464 19116 14516 19168
rect 15108 19116 15160 19168
rect 19156 19159 19208 19168
rect 19156 19125 19165 19159
rect 19165 19125 19199 19159
rect 19199 19125 19208 19159
rect 19156 19116 19208 19125
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 21824 19159 21876 19168
rect 21824 19125 21833 19159
rect 21833 19125 21867 19159
rect 21867 19125 21876 19159
rect 21824 19116 21876 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8484 18912 8536 18964
rect 9312 18912 9364 18964
rect 10876 18912 10928 18964
rect 14556 18912 14608 18964
rect 17500 18912 17552 18964
rect 10048 18844 10100 18896
rect 8300 18776 8352 18828
rect 10508 18776 10560 18828
rect 10968 18776 11020 18828
rect 12624 18776 12676 18828
rect 6552 18708 6604 18760
rect 10784 18708 10836 18760
rect 16396 18776 16448 18828
rect 19156 18776 19208 18828
rect 17500 18708 17552 18760
rect 23848 18819 23900 18828
rect 23848 18785 23857 18819
rect 23857 18785 23891 18819
rect 23891 18785 23900 18819
rect 23848 18776 23900 18785
rect 8300 18640 8352 18692
rect 8852 18640 8904 18692
rect 9404 18640 9456 18692
rect 8760 18572 8812 18624
rect 9220 18572 9272 18624
rect 10508 18640 10560 18692
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 11152 18640 11204 18692
rect 17684 18640 17736 18692
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22787 18751
rect 22787 18717 22796 18751
rect 22744 18708 22796 18717
rect 26792 18912 26844 18964
rect 24492 18640 24544 18692
rect 11520 18572 11572 18624
rect 12808 18572 12860 18624
rect 13268 18572 13320 18624
rect 14188 18572 14240 18624
rect 14280 18615 14332 18624
rect 14280 18581 14289 18615
rect 14289 18581 14323 18615
rect 14323 18581 14332 18615
rect 14280 18572 14332 18581
rect 17224 18572 17276 18624
rect 17500 18572 17552 18624
rect 20904 18572 20956 18624
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 24676 18615 24728 18624
rect 24676 18581 24685 18615
rect 24685 18581 24719 18615
rect 24719 18581 24728 18615
rect 24676 18572 24728 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 6552 18368 6604 18420
rect 9128 18368 9180 18420
rect 8208 18300 8260 18352
rect 10324 18368 10376 18420
rect 14188 18368 14240 18420
rect 11244 18300 11296 18352
rect 9496 18275 9548 18284
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 9588 18232 9640 18284
rect 7748 18207 7800 18216
rect 7748 18173 7757 18207
rect 7757 18173 7791 18207
rect 7791 18173 7800 18207
rect 7748 18164 7800 18173
rect 9680 18164 9732 18216
rect 7564 18028 7616 18080
rect 11336 18232 11388 18284
rect 12072 18300 12124 18352
rect 13360 18300 13412 18352
rect 11612 18232 11664 18284
rect 16580 18368 16632 18420
rect 25872 18368 25924 18420
rect 24860 18300 24912 18352
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 11244 18207 11296 18216
rect 11244 18173 11253 18207
rect 11253 18173 11287 18207
rect 11287 18173 11296 18207
rect 11244 18164 11296 18173
rect 11888 18164 11940 18216
rect 13452 18164 13504 18216
rect 16764 18164 16816 18216
rect 15016 18096 15068 18148
rect 16948 18028 17000 18080
rect 18328 18028 18380 18080
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 23480 18232 23532 18284
rect 24584 18207 24636 18216
rect 24584 18173 24593 18207
rect 24593 18173 24627 18207
rect 24627 18173 24636 18207
rect 24584 18164 24636 18173
rect 19156 18028 19208 18080
rect 21088 18071 21140 18080
rect 21088 18037 21097 18071
rect 21097 18037 21131 18071
rect 21131 18037 21140 18071
rect 21088 18028 21140 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9680 17824 9732 17876
rect 11244 17824 11296 17876
rect 14004 17824 14056 17876
rect 17868 17824 17920 17876
rect 7840 17688 7892 17740
rect 9496 17688 9548 17740
rect 10140 17688 10192 17740
rect 13452 17756 13504 17808
rect 13820 17756 13872 17808
rect 16672 17756 16724 17808
rect 23204 17756 23256 17808
rect 12532 17688 12584 17740
rect 17316 17688 17368 17740
rect 17684 17688 17736 17740
rect 18328 17688 18380 17740
rect 24860 17824 24912 17876
rect 26148 17756 26200 17808
rect 7656 17552 7708 17604
rect 7380 17527 7432 17536
rect 7380 17493 7389 17527
rect 7389 17493 7423 17527
rect 7423 17493 7432 17527
rect 7380 17484 7432 17493
rect 9404 17484 9456 17536
rect 11520 17620 11572 17672
rect 11888 17620 11940 17672
rect 14280 17620 14332 17672
rect 16764 17620 16816 17672
rect 17592 17620 17644 17672
rect 19432 17620 19484 17672
rect 11336 17552 11388 17604
rect 11980 17552 12032 17604
rect 10232 17484 10284 17536
rect 12072 17484 12124 17536
rect 14188 17552 14240 17604
rect 16304 17552 16356 17604
rect 13176 17484 13228 17536
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 17132 17484 17184 17536
rect 17776 17484 17828 17536
rect 18420 17484 18472 17536
rect 19248 17552 19300 17604
rect 21180 17620 21232 17672
rect 21916 17663 21968 17672
rect 21916 17629 21925 17663
rect 21925 17629 21959 17663
rect 21959 17629 21968 17663
rect 21916 17620 21968 17629
rect 22192 17620 22244 17672
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 23664 17620 23716 17672
rect 20720 17484 20772 17536
rect 24400 17552 24452 17604
rect 22560 17484 22612 17536
rect 24768 17484 24820 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 7380 17280 7432 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11060 17280 11112 17332
rect 9496 17212 9548 17264
rect 11336 17280 11388 17332
rect 11612 17323 11664 17332
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 12256 17280 12308 17332
rect 13176 17323 13228 17332
rect 13176 17289 13185 17323
rect 13185 17289 13219 17323
rect 13219 17289 13228 17323
rect 13176 17280 13228 17289
rect 15384 17280 15436 17332
rect 15752 17280 15804 17332
rect 17316 17280 17368 17332
rect 20168 17280 20220 17332
rect 22192 17280 22244 17332
rect 24124 17280 24176 17332
rect 15936 17212 15988 17264
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 8944 17144 8996 17196
rect 16856 17144 16908 17196
rect 17868 17212 17920 17264
rect 18512 17212 18564 17264
rect 18788 17212 18840 17264
rect 20996 17212 21048 17264
rect 21824 17212 21876 17264
rect 22284 17212 22336 17264
rect 23756 17255 23808 17264
rect 23756 17221 23765 17255
rect 23765 17221 23799 17255
rect 23799 17221 23808 17255
rect 23756 17212 23808 17221
rect 24032 17212 24084 17264
rect 8392 17076 8444 17128
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 12716 17076 12768 17128
rect 11520 17008 11572 17060
rect 12072 17051 12124 17060
rect 12072 17017 12081 17051
rect 12081 17017 12115 17051
rect 12115 17017 12124 17051
rect 12072 17008 12124 17017
rect 13636 17076 13688 17128
rect 14556 17119 14608 17128
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 14832 17076 14884 17128
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 20444 17008 20496 17060
rect 11796 16940 11848 16992
rect 16212 16940 16264 16992
rect 17592 16940 17644 16992
rect 22376 16940 22428 16992
rect 23204 16940 23256 16992
rect 23940 16940 23992 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 8392 16736 8444 16788
rect 11244 16711 11296 16720
rect 11244 16677 11253 16711
rect 11253 16677 11287 16711
rect 11287 16677 11296 16711
rect 11244 16668 11296 16677
rect 13268 16736 13320 16788
rect 14464 16736 14516 16788
rect 15752 16736 15804 16788
rect 12532 16600 12584 16652
rect 13176 16600 13228 16652
rect 13544 16643 13596 16652
rect 13544 16609 13553 16643
rect 13553 16609 13587 16643
rect 13587 16609 13596 16643
rect 13544 16600 13596 16609
rect 10416 16464 10468 16516
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 10600 16439 10652 16448
rect 9864 16396 9916 16405
rect 10600 16405 10609 16439
rect 10609 16405 10643 16439
rect 10643 16405 10652 16439
rect 10600 16396 10652 16405
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 16856 16600 16908 16652
rect 18604 16600 18656 16652
rect 15660 16532 15712 16584
rect 21272 16736 21324 16788
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 22744 16736 22796 16788
rect 23664 16736 23716 16788
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 20628 16600 20680 16652
rect 22284 16532 22336 16584
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 11796 16396 11848 16405
rect 14188 16439 14240 16448
rect 14188 16405 14197 16439
rect 14197 16405 14231 16439
rect 14231 16405 14240 16439
rect 14188 16396 14240 16405
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 16672 16464 16724 16516
rect 19340 16464 19392 16516
rect 16120 16396 16172 16448
rect 16488 16439 16540 16448
rect 16488 16405 16497 16439
rect 16497 16405 16531 16439
rect 16531 16405 16540 16439
rect 16488 16396 16540 16405
rect 16856 16439 16908 16448
rect 16856 16405 16865 16439
rect 16865 16405 16899 16439
rect 16899 16405 16908 16439
rect 16856 16396 16908 16405
rect 17316 16396 17368 16448
rect 19524 16396 19576 16448
rect 20996 16464 21048 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 13268 16192 13320 16244
rect 14188 16192 14240 16244
rect 14832 16192 14884 16244
rect 14924 16192 14976 16244
rect 16672 16192 16724 16244
rect 8300 16124 8352 16176
rect 8576 16124 8628 16176
rect 11336 16124 11388 16176
rect 13820 16124 13872 16176
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 14004 16056 14056 16108
rect 14740 16056 14792 16108
rect 17316 16167 17368 16176
rect 17316 16133 17325 16167
rect 17325 16133 17359 16167
rect 17359 16133 17368 16167
rect 17316 16124 17368 16133
rect 17960 16056 18012 16108
rect 18880 16124 18932 16176
rect 19340 16124 19392 16176
rect 19984 16192 20036 16244
rect 20260 16192 20312 16244
rect 20352 16124 20404 16176
rect 19984 16056 20036 16108
rect 23572 16192 23624 16244
rect 22284 16167 22336 16176
rect 22284 16133 22293 16167
rect 22293 16133 22327 16167
rect 22327 16133 22336 16167
rect 22284 16124 22336 16133
rect 22744 16124 22796 16176
rect 23848 16056 23900 16108
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 8668 15920 8720 15972
rect 11888 15920 11940 15972
rect 13636 15988 13688 16040
rect 13452 15920 13504 15972
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8576 15895 8628 15904
rect 8576 15861 8585 15895
rect 8585 15861 8619 15895
rect 8619 15861 8628 15895
rect 8576 15852 8628 15861
rect 13176 15852 13228 15904
rect 16580 15920 16632 15972
rect 22744 15988 22796 16040
rect 24032 16031 24084 16040
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 24584 15988 24636 16040
rect 16120 15852 16172 15904
rect 17224 15895 17276 15904
rect 17224 15861 17233 15895
rect 17233 15861 17267 15895
rect 17267 15861 17276 15895
rect 17224 15852 17276 15861
rect 19248 15852 19300 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 9036 15648 9088 15700
rect 11704 15648 11756 15700
rect 12624 15648 12676 15700
rect 14464 15648 14516 15700
rect 16396 15691 16448 15700
rect 16396 15657 16405 15691
rect 16405 15657 16439 15691
rect 16439 15657 16448 15691
rect 16396 15648 16448 15657
rect 11980 15580 12032 15632
rect 13452 15580 13504 15632
rect 15016 15580 15068 15632
rect 17316 15648 17368 15700
rect 18512 15648 18564 15700
rect 21456 15648 21508 15700
rect 24952 15648 25004 15700
rect 22744 15580 22796 15632
rect 24124 15580 24176 15632
rect 10692 15512 10744 15564
rect 11888 15512 11940 15564
rect 18604 15512 18656 15564
rect 20260 15512 20312 15564
rect 20720 15512 20772 15564
rect 6552 15444 6604 15496
rect 6828 15444 6880 15496
rect 9496 15444 9548 15496
rect 12256 15444 12308 15496
rect 22100 15512 22152 15564
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 23664 15512 23716 15564
rect 24768 15555 24820 15564
rect 24768 15521 24777 15555
rect 24777 15521 24811 15555
rect 24811 15521 24820 15555
rect 24768 15512 24820 15521
rect 12624 15376 12676 15428
rect 9404 15308 9456 15360
rect 12072 15351 12124 15360
rect 12072 15317 12081 15351
rect 12081 15317 12115 15351
rect 12115 15317 12124 15351
rect 12072 15308 12124 15317
rect 13728 15308 13780 15360
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 15936 15351 15988 15360
rect 15936 15317 15945 15351
rect 15945 15317 15979 15351
rect 15979 15317 15988 15351
rect 15936 15308 15988 15317
rect 16856 15308 16908 15360
rect 18328 15376 18380 15428
rect 19616 15376 19668 15428
rect 21272 15376 21324 15428
rect 22192 15376 22244 15428
rect 23756 15419 23808 15428
rect 23756 15385 23765 15419
rect 23765 15385 23799 15419
rect 23799 15385 23808 15419
rect 23756 15376 23808 15385
rect 19064 15308 19116 15360
rect 19800 15308 19852 15360
rect 20536 15308 20588 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 9956 15104 10008 15156
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 12256 15104 12308 15156
rect 14280 15104 14332 15156
rect 8668 15036 8720 15088
rect 15936 15147 15988 15156
rect 15936 15113 15945 15147
rect 15945 15113 15979 15147
rect 15979 15113 15988 15147
rect 15936 15104 15988 15113
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 17408 15104 17460 15156
rect 19892 15147 19944 15156
rect 19892 15113 19901 15147
rect 19901 15113 19935 15147
rect 19935 15113 19944 15147
rect 19892 15104 19944 15113
rect 21824 15104 21876 15156
rect 6828 14900 6880 14952
rect 8300 14900 8352 14952
rect 9312 14900 9364 14952
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11612 14968 11664 15020
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 12440 14900 12492 14952
rect 17040 15036 17092 15088
rect 20076 15036 20128 15088
rect 15200 14968 15252 15020
rect 14556 14900 14608 14952
rect 16948 14968 17000 15020
rect 18880 14968 18932 15020
rect 22836 15036 22888 15088
rect 23296 15079 23348 15088
rect 23296 15045 23305 15079
rect 23305 15045 23339 15079
rect 23339 15045 23348 15079
rect 23296 15036 23348 15045
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 12532 14807 12584 14816
rect 12532 14773 12541 14807
rect 12541 14773 12575 14807
rect 12575 14773 12584 14807
rect 12532 14764 12584 14773
rect 15476 14764 15528 14816
rect 19800 14943 19852 14952
rect 19800 14909 19809 14943
rect 19809 14909 19843 14943
rect 19843 14909 19852 14943
rect 19800 14900 19852 14909
rect 18604 14875 18656 14884
rect 18604 14841 18613 14875
rect 18613 14841 18647 14875
rect 18647 14841 18656 14875
rect 18604 14832 18656 14841
rect 19064 14832 19116 14884
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 22836 14832 22888 14884
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 7840 14560 7892 14612
rect 12808 14560 12860 14612
rect 20720 14560 20772 14612
rect 24308 14560 24360 14612
rect 15384 14535 15436 14544
rect 15384 14501 15393 14535
rect 15393 14501 15427 14535
rect 15427 14501 15436 14535
rect 15384 14492 15436 14501
rect 20812 14492 20864 14544
rect 7288 14424 7340 14476
rect 11244 14424 11296 14476
rect 12256 14424 12308 14476
rect 12992 14424 13044 14476
rect 9588 14356 9640 14408
rect 13820 14356 13872 14408
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15200 14424 15252 14476
rect 16028 14424 16080 14476
rect 19892 14356 19944 14408
rect 22008 14492 22060 14544
rect 23940 14492 23992 14544
rect 21732 14467 21784 14476
rect 21732 14433 21741 14467
rect 21741 14433 21775 14467
rect 21775 14433 21784 14467
rect 21732 14424 21784 14433
rect 24860 14424 24912 14476
rect 23296 14356 23348 14408
rect 24492 14356 24544 14408
rect 6828 14288 6880 14340
rect 10140 14288 10192 14340
rect 8668 14220 8720 14272
rect 11244 14220 11296 14272
rect 12164 14288 12216 14340
rect 14188 14288 14240 14340
rect 15384 14288 15436 14340
rect 19616 14288 19668 14340
rect 23388 14288 23440 14340
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 14372 14220 14424 14272
rect 15660 14220 15712 14272
rect 20168 14220 20220 14272
rect 20260 14263 20312 14272
rect 20260 14229 20269 14263
rect 20269 14229 20303 14263
rect 20303 14229 20312 14263
rect 20260 14220 20312 14229
rect 20444 14220 20496 14272
rect 23940 14220 23992 14272
rect 25136 14220 25188 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 9864 14016 9916 14068
rect 12992 14059 13044 14068
rect 12992 14025 13001 14059
rect 13001 14025 13035 14059
rect 13035 14025 13044 14059
rect 12992 14016 13044 14025
rect 14740 14016 14792 14068
rect 6828 13880 6880 13932
rect 8300 13948 8352 14000
rect 8668 13948 8720 14000
rect 11336 13948 11388 14000
rect 12256 13991 12308 14000
rect 12256 13957 12265 13991
rect 12265 13957 12299 13991
rect 12299 13957 12308 13991
rect 12256 13948 12308 13957
rect 16028 14016 16080 14068
rect 18788 14016 18840 14068
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 21180 14016 21232 14068
rect 22652 14016 22704 14068
rect 24032 14016 24084 14068
rect 19616 13991 19668 14000
rect 19616 13957 19625 13991
rect 19625 13957 19659 13991
rect 19659 13957 19668 13991
rect 19616 13948 19668 13957
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 9036 13812 9088 13864
rect 9588 13880 9640 13932
rect 10140 13812 10192 13864
rect 11888 13880 11940 13932
rect 12532 13880 12584 13932
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 12716 13812 12768 13864
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 16488 13812 16540 13864
rect 15200 13744 15252 13796
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 19064 13880 19116 13932
rect 20168 13923 20220 13932
rect 20168 13889 20177 13923
rect 20177 13889 20211 13923
rect 20211 13889 20220 13923
rect 20168 13880 20220 13889
rect 22468 13948 22520 14000
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 24216 13880 24268 13932
rect 24400 13880 24452 13932
rect 14096 13719 14148 13728
rect 14096 13685 14126 13719
rect 14126 13685 14148 13719
rect 14096 13676 14148 13685
rect 17316 13676 17368 13728
rect 17592 13676 17644 13728
rect 18512 13744 18564 13796
rect 21272 13812 21324 13864
rect 22192 13812 22244 13864
rect 23204 13812 23256 13864
rect 20996 13676 21048 13728
rect 22284 13676 22336 13728
rect 22652 13676 22704 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 7656 13472 7708 13524
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 14556 13472 14608 13524
rect 15660 13472 15712 13524
rect 15752 13472 15804 13524
rect 16672 13472 16724 13524
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 17592 13472 17644 13524
rect 24216 13472 24268 13524
rect 24492 13472 24544 13524
rect 13268 13404 13320 13456
rect 15568 13404 15620 13456
rect 21088 13447 21140 13456
rect 21088 13413 21097 13447
rect 21097 13413 21131 13447
rect 21131 13413 21140 13447
rect 21088 13404 21140 13413
rect 21180 13404 21232 13456
rect 7288 13336 7340 13388
rect 11520 13336 11572 13388
rect 13820 13336 13872 13388
rect 15292 13336 15344 13388
rect 15936 13336 15988 13388
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 9036 13268 9088 13320
rect 13912 13268 13964 13320
rect 14924 13268 14976 13320
rect 16120 13268 16172 13320
rect 9128 13200 9180 13252
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 11244 13200 11296 13252
rect 11796 13200 11848 13252
rect 12164 13200 12216 13252
rect 15476 13200 15528 13252
rect 20076 13336 20128 13388
rect 23388 13379 23440 13388
rect 23388 13345 23397 13379
rect 23397 13345 23431 13379
rect 23431 13345 23440 13379
rect 23388 13336 23440 13345
rect 17408 13268 17460 13320
rect 18328 13268 18380 13320
rect 17040 13200 17092 13252
rect 18512 13243 18564 13252
rect 18512 13209 18521 13243
rect 18521 13209 18555 13243
rect 18555 13209 18564 13243
rect 18512 13200 18564 13209
rect 12348 13132 12400 13184
rect 14924 13175 14976 13184
rect 14924 13141 14933 13175
rect 14933 13141 14967 13175
rect 14967 13141 14976 13175
rect 14924 13132 14976 13141
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 19340 13268 19392 13320
rect 21916 13311 21968 13320
rect 21916 13277 21925 13311
rect 21925 13277 21959 13311
rect 21959 13277 21968 13311
rect 21916 13268 21968 13277
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 24308 13200 24360 13252
rect 24400 13200 24452 13252
rect 22192 13132 22244 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 7564 12928 7616 12980
rect 9496 12928 9548 12980
rect 11704 12928 11756 12980
rect 12256 12928 12308 12980
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 14832 12928 14884 12980
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 17132 12971 17184 12980
rect 17132 12937 17141 12971
rect 17141 12937 17175 12971
rect 17175 12937 17184 12971
rect 17132 12928 17184 12937
rect 17592 12971 17644 12980
rect 17592 12937 17601 12971
rect 17601 12937 17635 12971
rect 17635 12937 17644 12971
rect 17592 12928 17644 12937
rect 6920 12860 6972 12912
rect 9864 12860 9916 12912
rect 7380 12792 7432 12844
rect 7840 12792 7892 12844
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 8944 12792 8996 12844
rect 11244 12860 11296 12912
rect 8484 12724 8536 12776
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 10048 12724 10100 12776
rect 13268 12792 13320 12844
rect 13636 12792 13688 12844
rect 15568 12860 15620 12912
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 19984 12928 20036 12980
rect 22008 12928 22060 12980
rect 22100 12928 22152 12980
rect 23480 12928 23532 12980
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12256 12724 12308 12776
rect 7012 12656 7064 12708
rect 9404 12656 9456 12708
rect 10784 12656 10836 12708
rect 12532 12656 12584 12708
rect 13820 12724 13872 12776
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 15292 12724 15344 12776
rect 15476 12724 15528 12776
rect 15384 12656 15436 12708
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 18328 12792 18380 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 22376 12860 22428 12912
rect 23296 12860 23348 12912
rect 24400 12928 24452 12980
rect 20628 12792 20680 12844
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 22100 12792 22152 12844
rect 22192 12792 22244 12844
rect 18788 12724 18840 12776
rect 20628 12656 20680 12708
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 11152 12588 11204 12640
rect 11796 12588 11848 12640
rect 12716 12588 12768 12640
rect 13452 12588 13504 12640
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 23388 12588 23440 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 10232 12427 10284 12436
rect 10232 12393 10241 12427
rect 10241 12393 10275 12427
rect 10275 12393 10284 12427
rect 10232 12384 10284 12393
rect 10508 12384 10560 12436
rect 11980 12384 12032 12436
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 12440 12316 12492 12368
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 13544 12384 13596 12436
rect 12716 12316 12768 12368
rect 14096 12384 14148 12436
rect 14832 12384 14884 12436
rect 7288 12180 7340 12232
rect 10968 12248 11020 12300
rect 12164 12248 12216 12300
rect 12532 12248 12584 12300
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 14004 12248 14056 12300
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 14832 12291 14884 12300
rect 14832 12257 14841 12291
rect 14841 12257 14875 12291
rect 14875 12257 14884 12291
rect 14832 12248 14884 12257
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 18788 12384 18840 12436
rect 19432 12384 19484 12436
rect 19892 12384 19944 12436
rect 21364 12384 21416 12436
rect 24124 12384 24176 12436
rect 15108 12316 15160 12368
rect 15476 12359 15528 12368
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 16028 12316 16080 12368
rect 19064 12316 19116 12368
rect 20260 12316 20312 12368
rect 20536 12316 20588 12368
rect 22560 12316 22612 12368
rect 22836 12316 22888 12368
rect 12532 12112 12584 12164
rect 18696 12248 18748 12300
rect 19156 12248 19208 12300
rect 19340 12180 19392 12232
rect 20720 12248 20772 12300
rect 21272 12248 21324 12300
rect 24860 12248 24912 12300
rect 22192 12223 22244 12232
rect 22192 12189 22201 12223
rect 22201 12189 22235 12223
rect 22235 12189 22244 12223
rect 22192 12180 22244 12189
rect 22836 12180 22888 12232
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 24124 12180 24176 12232
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 12716 12044 12768 12096
rect 13912 12044 13964 12096
rect 16948 12112 17000 12164
rect 17408 12155 17460 12164
rect 17408 12121 17417 12155
rect 17417 12121 17451 12155
rect 17451 12121 17460 12155
rect 17408 12112 17460 12121
rect 19892 12112 19944 12164
rect 21364 12112 21416 12164
rect 15384 12044 15436 12096
rect 15844 12044 15896 12096
rect 18420 12044 18472 12096
rect 20352 12044 20404 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 8668 11840 8720 11892
rect 9588 11840 9640 11892
rect 9680 11840 9732 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 11336 11840 11388 11892
rect 11980 11840 12032 11892
rect 12808 11840 12860 11892
rect 13084 11840 13136 11892
rect 13544 11840 13596 11892
rect 14464 11840 14516 11892
rect 14740 11840 14792 11892
rect 15660 11840 15712 11892
rect 17500 11840 17552 11892
rect 17868 11840 17920 11892
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 18880 11840 18932 11892
rect 9128 11636 9180 11688
rect 3976 11500 4028 11552
rect 14372 11772 14424 11824
rect 11060 11636 11112 11688
rect 11888 11636 11940 11688
rect 10232 11568 10284 11620
rect 9680 11500 9732 11552
rect 9864 11500 9916 11552
rect 11980 11500 12032 11552
rect 14556 11704 14608 11756
rect 16488 11772 16540 11824
rect 16672 11772 16724 11824
rect 16764 11772 16816 11824
rect 17592 11772 17644 11824
rect 12808 11636 12860 11688
rect 13084 11611 13136 11620
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 16488 11636 16540 11688
rect 19800 11772 19852 11824
rect 20352 11840 20404 11892
rect 20720 11840 20772 11892
rect 21456 11883 21508 11892
rect 21456 11849 21465 11883
rect 21465 11849 21499 11883
rect 21499 11849 21508 11883
rect 21456 11840 21508 11849
rect 20076 11815 20128 11824
rect 20076 11781 20085 11815
rect 20085 11781 20119 11815
rect 20119 11781 20128 11815
rect 20076 11772 20128 11781
rect 25964 11772 26016 11824
rect 19432 11704 19484 11756
rect 20352 11704 20404 11756
rect 20904 11704 20956 11756
rect 24400 11704 24452 11756
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 19984 11636 20036 11688
rect 14648 11500 14700 11552
rect 15292 11500 15344 11552
rect 16396 11500 16448 11552
rect 21456 11568 21508 11620
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 24860 11568 24912 11620
rect 18604 11500 18656 11552
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 20168 11543 20220 11552
rect 20168 11509 20177 11543
rect 20177 11509 20211 11543
rect 20211 11509 20220 11543
rect 20168 11500 20220 11509
rect 20260 11500 20312 11552
rect 21824 11500 21876 11552
rect 23296 11500 23348 11552
rect 25780 11500 25832 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 12716 11296 12768 11348
rect 12900 11296 12952 11348
rect 12992 11296 13044 11348
rect 15200 11296 15252 11348
rect 16304 11296 16356 11348
rect 10600 11228 10652 11280
rect 12624 11228 12676 11280
rect 10416 11160 10468 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 11060 11092 11112 11144
rect 13544 11160 13596 11212
rect 13912 11228 13964 11280
rect 14464 11228 14516 11280
rect 16488 11228 16540 11280
rect 17040 11228 17092 11280
rect 17316 11228 17368 11280
rect 17868 11339 17920 11348
rect 17868 11305 17877 11339
rect 17877 11305 17911 11339
rect 17911 11305 17920 11339
rect 17868 11296 17920 11305
rect 20260 11296 20312 11348
rect 20444 11296 20496 11348
rect 20720 11296 20772 11348
rect 23296 11296 23348 11348
rect 24032 11296 24084 11348
rect 20628 11228 20680 11280
rect 22744 11228 22796 11280
rect 14096 11160 14148 11212
rect 15936 11160 15988 11212
rect 17408 11160 17460 11212
rect 19340 11160 19392 11212
rect 22652 11160 22704 11212
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 14832 11092 14884 11144
rect 18788 11092 18840 11144
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20720 11092 20772 11144
rect 21456 11092 21508 11144
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 10416 11024 10468 11076
rect 12532 11024 12584 11076
rect 11796 10999 11848 11008
rect 11796 10965 11805 10999
rect 11805 10965 11839 10999
rect 11839 10965 11848 10999
rect 11796 10956 11848 10965
rect 12716 11024 12768 11076
rect 14464 11024 14516 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 16672 11024 16724 11076
rect 17316 11024 17368 11076
rect 20812 11067 20864 11076
rect 20812 11033 20821 11067
rect 20821 11033 20855 11067
rect 20855 11033 20864 11067
rect 20812 11024 20864 11033
rect 12992 10999 13044 11008
rect 12992 10965 13001 10999
rect 13001 10965 13035 10999
rect 13035 10965 13044 10999
rect 12992 10956 13044 10965
rect 15016 10956 15068 11008
rect 19800 10956 19852 11008
rect 19984 10956 20036 11008
rect 21456 10956 21508 11008
rect 21732 10999 21784 11008
rect 21732 10965 21741 10999
rect 21741 10965 21775 10999
rect 21775 10965 21784 10999
rect 21732 10956 21784 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 10048 10752 10100 10804
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 14188 10752 14240 10804
rect 7104 10412 7156 10464
rect 9864 10684 9916 10736
rect 10416 10684 10468 10736
rect 11888 10684 11940 10736
rect 15476 10752 15528 10804
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 16304 10752 16356 10804
rect 19984 10752 20036 10804
rect 22192 10752 22244 10804
rect 14188 10659 14240 10668
rect 14188 10625 14197 10659
rect 14197 10625 14231 10659
rect 14231 10625 14240 10659
rect 14188 10616 14240 10625
rect 8484 10548 8536 10600
rect 11796 10548 11848 10600
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 10600 10480 10652 10532
rect 12900 10548 12952 10600
rect 13728 10548 13780 10600
rect 13912 10548 13964 10600
rect 9128 10412 9180 10464
rect 9588 10412 9640 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10968 10455 11020 10464
rect 10416 10412 10468 10421
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 18328 10684 18380 10736
rect 15476 10616 15528 10668
rect 16856 10659 16908 10668
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 17776 10616 17828 10668
rect 15292 10548 15344 10600
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 19616 10684 19668 10736
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 15568 10412 15620 10464
rect 17500 10523 17552 10532
rect 17500 10489 17509 10523
rect 17509 10489 17543 10523
rect 17543 10489 17552 10523
rect 17500 10480 17552 10489
rect 19984 10616 20036 10668
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 22284 10616 22336 10668
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 20444 10548 20496 10600
rect 20628 10548 20680 10600
rect 21272 10591 21324 10600
rect 21272 10557 21281 10591
rect 21281 10557 21315 10591
rect 21315 10557 21324 10591
rect 21272 10548 21324 10557
rect 21456 10548 21508 10600
rect 24124 10752 24176 10804
rect 23388 10727 23440 10736
rect 23388 10693 23397 10727
rect 23397 10693 23431 10727
rect 23431 10693 23440 10727
rect 23388 10684 23440 10693
rect 25320 10684 25372 10736
rect 22836 10548 22888 10600
rect 18788 10412 18840 10464
rect 21640 10480 21692 10532
rect 22100 10480 22152 10532
rect 22008 10455 22060 10464
rect 22008 10421 22017 10455
rect 22017 10421 22051 10455
rect 22051 10421 22060 10455
rect 22008 10412 22060 10421
rect 22468 10455 22520 10464
rect 22468 10421 22477 10455
rect 22477 10421 22511 10455
rect 22511 10421 22520 10455
rect 22468 10412 22520 10421
rect 22744 10455 22796 10464
rect 22744 10421 22753 10455
rect 22753 10421 22787 10455
rect 22787 10421 22796 10455
rect 22744 10412 22796 10421
rect 23480 10412 23532 10464
rect 24124 10412 24176 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 9588 10072 9640 10124
rect 10140 10072 10192 10124
rect 13728 10208 13780 10260
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 16028 10208 16080 10260
rect 19984 10208 20036 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12348 10072 12400 10124
rect 13544 10072 13596 10124
rect 11888 10004 11940 10056
rect 9312 9936 9364 9988
rect 10968 9936 11020 9988
rect 11612 9936 11664 9988
rect 13728 9936 13780 9988
rect 14188 10140 14240 10192
rect 16580 10140 16632 10192
rect 20536 10140 20588 10192
rect 14464 10072 14516 10124
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 14740 10004 14792 10056
rect 17684 10004 17736 10056
rect 17868 9936 17920 9988
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 19340 10072 19392 10124
rect 20904 10072 20956 10124
rect 21364 10072 21416 10124
rect 21548 10072 21600 10124
rect 24124 10072 24176 10124
rect 18972 10004 19024 10056
rect 22560 10004 22612 10056
rect 20260 9936 20312 9988
rect 21364 9936 21416 9988
rect 22192 9936 22244 9988
rect 25044 9936 25096 9988
rect 12808 9868 12860 9920
rect 13452 9868 13504 9920
rect 15476 9868 15528 9920
rect 15568 9868 15620 9920
rect 16028 9868 16080 9920
rect 16396 9868 16448 9920
rect 16764 9868 16816 9920
rect 18236 9868 18288 9920
rect 19524 9911 19576 9920
rect 19524 9877 19533 9911
rect 19533 9877 19567 9911
rect 19567 9877 19576 9911
rect 19524 9868 19576 9877
rect 19800 9868 19852 9920
rect 19984 9911 20036 9920
rect 19984 9877 19993 9911
rect 19993 9877 20027 9911
rect 20027 9877 20036 9911
rect 19984 9868 20036 9877
rect 21640 9868 21692 9920
rect 22376 9868 22428 9920
rect 24584 9868 24636 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 7104 9664 7156 9716
rect 12348 9664 12400 9716
rect 15292 9664 15344 9716
rect 15476 9664 15528 9716
rect 17408 9664 17460 9716
rect 18972 9664 19024 9716
rect 3884 9596 3936 9648
rect 8852 9596 8904 9648
rect 11612 9596 11664 9648
rect 16120 9596 16172 9648
rect 16304 9596 16356 9648
rect 16672 9596 16724 9648
rect 16948 9596 17000 9648
rect 15384 9528 15436 9580
rect 10692 9460 10744 9512
rect 11520 9460 11572 9512
rect 12716 9460 12768 9512
rect 13820 9460 13872 9512
rect 14004 9460 14056 9512
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 13728 9392 13780 9444
rect 14832 9392 14884 9444
rect 17316 9528 17368 9580
rect 15660 9460 15712 9512
rect 15844 9460 15896 9512
rect 16028 9460 16080 9512
rect 18696 9596 18748 9648
rect 19800 9596 19852 9648
rect 20904 9664 20956 9716
rect 21088 9664 21140 9716
rect 20720 9596 20772 9648
rect 21456 9596 21508 9648
rect 21548 9596 21600 9648
rect 22744 9596 22796 9648
rect 23388 9664 23440 9716
rect 25320 9707 25372 9716
rect 25320 9673 25329 9707
rect 25329 9673 25363 9707
rect 25363 9673 25372 9707
rect 25320 9664 25372 9673
rect 23480 9596 23532 9648
rect 24124 9639 24176 9648
rect 24124 9605 24133 9639
rect 24133 9605 24167 9639
rect 24167 9605 24176 9639
rect 24124 9596 24176 9605
rect 19248 9528 19300 9580
rect 22560 9528 22612 9580
rect 24952 9528 25004 9580
rect 11520 9324 11572 9376
rect 14372 9324 14424 9376
rect 16580 9392 16632 9444
rect 17040 9392 17092 9444
rect 22652 9503 22704 9512
rect 22652 9469 22661 9503
rect 22661 9469 22695 9503
rect 22695 9469 22704 9503
rect 22652 9460 22704 9469
rect 19800 9392 19852 9444
rect 22100 9392 22152 9444
rect 22836 9392 22888 9444
rect 16672 9324 16724 9376
rect 17408 9324 17460 9376
rect 21364 9324 21416 9376
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 12348 9120 12400 9172
rect 12624 9120 12676 9172
rect 12808 9120 12860 9172
rect 15752 9120 15804 9172
rect 16672 9120 16724 9172
rect 17960 9120 18012 9172
rect 19340 9120 19392 9172
rect 12440 9052 12492 9104
rect 14004 9052 14056 9104
rect 15660 9052 15712 9104
rect 17040 9052 17092 9104
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14464 8984 14516 9036
rect 16304 8984 16356 9036
rect 17684 9027 17736 9036
rect 17684 8993 17693 9027
rect 17693 8993 17727 9027
rect 17727 8993 17736 9027
rect 17684 8984 17736 8993
rect 9312 8780 9364 8832
rect 10692 8848 10744 8900
rect 12624 8916 12676 8968
rect 16028 8916 16080 8968
rect 19984 9052 20036 9104
rect 17960 8984 18012 9036
rect 19064 8984 19116 9036
rect 20996 8984 21048 9036
rect 22100 8984 22152 9036
rect 19156 8916 19208 8968
rect 21456 8916 21508 8968
rect 13544 8848 13596 8900
rect 13820 8848 13872 8900
rect 14832 8848 14884 8900
rect 11520 8780 11572 8832
rect 14188 8780 14240 8832
rect 14556 8780 14608 8832
rect 15292 8780 15344 8832
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 15568 8780 15620 8832
rect 17408 8780 17460 8832
rect 17868 8848 17920 8900
rect 18420 8848 18472 8900
rect 19524 8848 19576 8900
rect 19800 8848 19852 8900
rect 20352 8780 20404 8832
rect 21180 8848 21232 8900
rect 24216 8916 24268 8968
rect 24952 8848 25004 8900
rect 21272 8780 21324 8832
rect 22192 8780 22244 8832
rect 23388 8780 23440 8832
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 13360 8576 13412 8628
rect 14096 8576 14148 8628
rect 21180 8576 21232 8628
rect 14464 8551 14516 8560
rect 14464 8517 14473 8551
rect 14473 8517 14507 8551
rect 14507 8517 14516 8551
rect 14464 8508 14516 8517
rect 14372 8440 14424 8492
rect 15016 8440 15068 8492
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 13912 8372 13964 8424
rect 17316 8440 17368 8492
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 15660 8415 15712 8424
rect 15660 8381 15669 8415
rect 15669 8381 15703 8415
rect 15703 8381 15712 8415
rect 15660 8372 15712 8381
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 17040 8415 17092 8424
rect 17040 8381 17049 8415
rect 17049 8381 17083 8415
rect 17083 8381 17092 8415
rect 17040 8372 17092 8381
rect 14832 8304 14884 8356
rect 15384 8304 15436 8356
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 20444 8415 20496 8424
rect 20444 8381 20453 8415
rect 20453 8381 20487 8415
rect 20487 8381 20496 8415
rect 20444 8372 20496 8381
rect 20628 8304 20680 8356
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 22192 8440 22244 8492
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 22468 8372 22520 8424
rect 21548 8304 21600 8356
rect 21824 8304 21876 8356
rect 24124 8304 24176 8356
rect 16212 8236 16264 8288
rect 22008 8236 22060 8288
rect 24492 8236 24544 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 10324 8032 10376 8084
rect 14096 8032 14148 8084
rect 14188 8032 14240 8084
rect 11796 8007 11848 8016
rect 11796 7973 11805 8007
rect 11805 7973 11839 8007
rect 11839 7973 11848 8007
rect 11796 7964 11848 7973
rect 12716 7964 12768 8016
rect 11888 7896 11940 7948
rect 17776 7964 17828 8016
rect 11704 7828 11756 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 15200 7896 15252 7948
rect 15844 7896 15896 7948
rect 17684 7896 17736 7948
rect 25320 8032 25372 8084
rect 23480 7964 23532 8016
rect 24032 7964 24084 8016
rect 16120 7828 16172 7880
rect 8576 7760 8628 7812
rect 17224 7828 17276 7880
rect 20076 7828 20128 7880
rect 11336 7735 11388 7744
rect 11336 7701 11345 7735
rect 11345 7701 11379 7735
rect 11379 7701 11388 7735
rect 11336 7692 11388 7701
rect 12624 7692 12676 7744
rect 16304 7803 16356 7812
rect 16304 7769 16313 7803
rect 16313 7769 16347 7803
rect 16347 7769 16356 7803
rect 16304 7760 16356 7769
rect 16396 7760 16448 7812
rect 21088 7760 21140 7812
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 15292 7692 15344 7744
rect 15844 7692 15896 7744
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 19340 7692 19392 7744
rect 19800 7692 19852 7744
rect 22836 7896 22888 7948
rect 21824 7828 21876 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 23388 7828 23440 7880
rect 22560 7692 22612 7744
rect 23664 7760 23716 7812
rect 24676 7692 24728 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 16856 7488 16908 7540
rect 18328 7488 18380 7540
rect 9588 7420 9640 7472
rect 11520 7420 11572 7472
rect 14464 7420 14516 7472
rect 16488 7420 16540 7472
rect 16948 7420 17000 7472
rect 17868 7420 17920 7472
rect 12072 7352 12124 7404
rect 13820 7352 13872 7404
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 12532 7327 12584 7336
rect 12532 7293 12541 7327
rect 12541 7293 12575 7327
rect 12575 7293 12584 7327
rect 12532 7284 12584 7293
rect 15108 7284 15160 7336
rect 11520 7216 11572 7268
rect 11888 7216 11940 7268
rect 15936 7284 15988 7336
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 11428 7148 11480 7200
rect 13544 7148 13596 7200
rect 17408 7216 17460 7268
rect 16580 7148 16632 7200
rect 16948 7148 17000 7200
rect 18696 7488 18748 7540
rect 19800 7488 19852 7540
rect 20628 7488 20680 7540
rect 20536 7420 20588 7472
rect 22100 7420 22152 7472
rect 23388 7420 23440 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 23848 7352 23900 7404
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 18604 7284 18656 7336
rect 21272 7327 21324 7336
rect 21272 7293 21281 7327
rect 21281 7293 21315 7327
rect 21315 7293 21324 7327
rect 21272 7284 21324 7293
rect 24860 7284 24912 7336
rect 21180 7216 21232 7268
rect 20904 7148 20956 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 17408 6944 17460 6996
rect 18696 6944 18748 6996
rect 13360 6876 13412 6928
rect 13636 6876 13688 6928
rect 16304 6876 16356 6928
rect 12716 6808 12768 6860
rect 10692 6740 10744 6792
rect 11060 6715 11112 6724
rect 11060 6681 11069 6715
rect 11069 6681 11103 6715
rect 11103 6681 11112 6715
rect 11060 6672 11112 6681
rect 4068 6604 4120 6656
rect 9772 6604 9824 6656
rect 11520 6672 11572 6724
rect 14464 6808 14516 6860
rect 15936 6808 15988 6860
rect 19800 6876 19852 6928
rect 21456 6876 21508 6928
rect 22836 6876 22888 6928
rect 23480 6876 23532 6928
rect 13728 6740 13780 6792
rect 21640 6808 21692 6860
rect 23296 6808 23348 6860
rect 25044 6851 25096 6860
rect 25044 6817 25053 6851
rect 25053 6817 25087 6851
rect 25087 6817 25096 6851
rect 25044 6808 25096 6817
rect 14648 6672 14700 6724
rect 13636 6604 13688 6656
rect 14372 6604 14424 6656
rect 16488 6672 16540 6724
rect 17040 6672 17092 6724
rect 17684 6672 17736 6724
rect 17868 6672 17920 6724
rect 21272 6740 21324 6792
rect 22008 6783 22060 6792
rect 22008 6749 22017 6783
rect 22017 6749 22051 6783
rect 22051 6749 22060 6783
rect 22008 6740 22060 6749
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 19156 6604 19208 6656
rect 20076 6604 20128 6656
rect 20996 6672 21048 6724
rect 21548 6672 21600 6724
rect 22376 6672 22428 6724
rect 24860 6672 24912 6724
rect 25228 6672 25280 6724
rect 20628 6604 20680 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 12808 6443 12860 6452
rect 12808 6409 12817 6443
rect 12817 6409 12851 6443
rect 12851 6409 12860 6443
rect 12808 6400 12860 6409
rect 17868 6400 17920 6452
rect 18972 6400 19024 6452
rect 20628 6400 20680 6452
rect 21640 6400 21692 6452
rect 11428 6332 11480 6384
rect 13820 6332 13872 6384
rect 6644 6264 6696 6316
rect 9312 6196 9364 6248
rect 6736 6128 6788 6180
rect 12164 6264 12216 6316
rect 11060 6196 11112 6248
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 14096 6196 14148 6248
rect 16120 6196 16172 6248
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 17776 6264 17828 6316
rect 19156 6332 19208 6384
rect 20260 6332 20312 6384
rect 21548 6332 21600 6384
rect 23388 6332 23440 6384
rect 24400 6400 24452 6452
rect 24676 6400 24728 6452
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 21456 6307 21508 6316
rect 21456 6273 21465 6307
rect 21465 6273 21499 6307
rect 21499 6273 21508 6307
rect 21456 6264 21508 6273
rect 23388 6196 23440 6248
rect 23480 6239 23532 6248
rect 23480 6205 23489 6239
rect 23489 6205 23523 6239
rect 23523 6205 23532 6239
rect 23480 6196 23532 6205
rect 24032 6239 24084 6248
rect 24032 6205 24041 6239
rect 24041 6205 24075 6239
rect 24075 6205 24084 6239
rect 24032 6196 24084 6205
rect 12532 6128 12584 6180
rect 14556 6128 14608 6180
rect 14648 6128 14700 6180
rect 14464 6060 14516 6112
rect 21732 6060 21784 6112
rect 24216 6103 24268 6112
rect 24216 6069 24225 6103
rect 24225 6069 24259 6103
rect 24259 6069 24268 6103
rect 24216 6060 24268 6069
rect 25228 6103 25280 6112
rect 25228 6069 25237 6103
rect 25237 6069 25271 6103
rect 25271 6069 25280 6103
rect 25228 6060 25280 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 13820 5856 13872 5908
rect 16856 5856 16908 5908
rect 11428 5788 11480 5840
rect 12992 5788 13044 5840
rect 14096 5788 14148 5840
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 17776 5856 17828 5908
rect 21456 5856 21508 5908
rect 23756 5856 23808 5908
rect 24308 5856 24360 5908
rect 10784 5720 10836 5772
rect 11060 5720 11112 5772
rect 12440 5720 12492 5772
rect 9588 5652 9640 5704
rect 11428 5652 11480 5704
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 13452 5652 13504 5704
rect 15384 5720 15436 5772
rect 19340 5720 19392 5772
rect 19708 5720 19760 5772
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 20812 5695 20864 5704
rect 20812 5661 20821 5695
rect 20821 5661 20855 5695
rect 20855 5661 20864 5695
rect 20812 5652 20864 5661
rect 22284 5652 22336 5704
rect 24216 5720 24268 5772
rect 23940 5652 23992 5704
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 14464 5627 14516 5636
rect 14464 5593 14473 5627
rect 14473 5593 14507 5627
rect 14507 5593 14516 5627
rect 14464 5584 14516 5593
rect 19340 5584 19392 5636
rect 20720 5584 20772 5636
rect 23756 5584 23808 5636
rect 12992 5516 13044 5568
rect 15292 5516 15344 5568
rect 16396 5516 16448 5568
rect 18328 5516 18380 5568
rect 22744 5516 22796 5568
rect 23296 5516 23348 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 11796 5244 11848 5296
rect 10968 5176 11020 5228
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 13544 5244 13596 5296
rect 14464 5244 14516 5296
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 10692 5040 10744 5092
rect 10600 4972 10652 5024
rect 15292 5244 15344 5296
rect 14924 5108 14976 5160
rect 16948 5176 17000 5228
rect 15752 5151 15804 5160
rect 15752 5117 15761 5151
rect 15761 5117 15795 5151
rect 15795 5117 15804 5151
rect 15752 5108 15804 5117
rect 15844 5108 15896 5160
rect 17040 5108 17092 5160
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 22744 5312 22796 5364
rect 19800 5244 19852 5296
rect 20260 5244 20312 5296
rect 21088 5244 21140 5296
rect 20536 5219 20588 5228
rect 20536 5185 20545 5219
rect 20545 5185 20579 5219
rect 20579 5185 20588 5219
rect 20536 5176 20588 5185
rect 21272 5244 21324 5296
rect 21456 5176 21508 5228
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 23756 5176 23808 5228
rect 18420 5108 18472 5160
rect 18604 5108 18656 5160
rect 21088 5108 21140 5160
rect 21272 5108 21324 5160
rect 23572 5108 23624 5160
rect 13912 4972 13964 5024
rect 14188 4972 14240 5024
rect 17408 4972 17460 5024
rect 17684 4972 17736 5024
rect 22652 4972 22704 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 14280 4768 14332 4820
rect 9588 4632 9640 4684
rect 10324 4675 10376 4684
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 11428 4700 11480 4752
rect 16856 4811 16908 4820
rect 16856 4777 16865 4811
rect 16865 4777 16899 4811
rect 16899 4777 16908 4811
rect 16856 4768 16908 4777
rect 17040 4768 17092 4820
rect 23756 4768 23808 4820
rect 10968 4632 11020 4684
rect 18604 4700 18656 4752
rect 14924 4632 14976 4684
rect 15936 4632 15988 4684
rect 20536 4632 20588 4684
rect 9680 4496 9732 4548
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 19616 4564 19668 4616
rect 21732 4607 21784 4616
rect 21732 4573 21741 4607
rect 21741 4573 21775 4607
rect 21775 4573 21784 4607
rect 21732 4564 21784 4573
rect 21824 4564 21876 4616
rect 15292 4496 15344 4548
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 16396 4496 16448 4548
rect 17316 4496 17368 4548
rect 20536 4496 20588 4548
rect 21640 4496 21692 4548
rect 22376 4496 22428 4548
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 11612 4428 11664 4480
rect 17224 4428 17276 4480
rect 21088 4428 21140 4480
rect 21364 4428 21416 4480
rect 23756 4539 23808 4548
rect 23756 4505 23765 4539
rect 23765 4505 23799 4539
rect 23799 4505 23808 4539
rect 23756 4496 23808 4505
rect 23664 4471 23716 4480
rect 23664 4437 23673 4471
rect 23673 4437 23707 4471
rect 23707 4437 23716 4471
rect 23664 4428 23716 4437
rect 24308 4428 24360 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 1492 4088 1544 4140
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 15476 4224 15528 4276
rect 17868 4224 17920 4276
rect 22008 4224 22060 4276
rect 4068 4088 4120 4140
rect 5908 4088 5960 4140
rect 14188 4199 14240 4208
rect 14188 4165 14197 4199
rect 14197 4165 14231 4199
rect 14231 4165 14240 4199
rect 14188 4156 14240 4165
rect 16396 4156 16448 4208
rect 19800 4156 19852 4208
rect 20536 4156 20588 4208
rect 8944 4088 8996 4140
rect 9220 4088 9272 4140
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 3700 3952 3752 4004
rect 7012 4020 7064 4072
rect 5908 3952 5960 4004
rect 6552 3952 6604 4004
rect 12440 4020 12492 4072
rect 12808 4020 12860 4072
rect 16028 4020 16080 4072
rect 16212 4020 16264 4072
rect 18512 4088 18564 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 21456 4156 21508 4208
rect 24216 4131 24268 4140
rect 24216 4097 24225 4131
rect 24225 4097 24259 4131
rect 24259 4097 24268 4131
rect 24216 4088 24268 4097
rect 24308 4088 24360 4140
rect 18328 4020 18380 4072
rect 18420 4020 18472 4072
rect 21088 4063 21140 4072
rect 21088 4029 21097 4063
rect 21097 4029 21131 4063
rect 21131 4029 21140 4063
rect 21088 4020 21140 4029
rect 2688 3884 2740 3936
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 4068 3884 4120 3936
rect 5264 3884 5316 3936
rect 5448 3884 5500 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 7196 3884 7248 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 11060 3884 11112 3936
rect 11888 3884 11940 3936
rect 15660 3952 15712 4004
rect 20260 3952 20312 4004
rect 21272 3952 21324 4004
rect 18880 3884 18932 3936
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 25228 3884 25280 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 1584 3680 1636 3732
rect 7840 3680 7892 3732
rect 8576 3723 8628 3732
rect 8576 3689 8585 3723
rect 8585 3689 8619 3723
rect 8619 3689 8628 3723
rect 8576 3680 8628 3689
rect 13820 3680 13872 3732
rect 19248 3680 19300 3732
rect 20352 3680 20404 3732
rect 22928 3680 22980 3732
rect 24216 3680 24268 3732
rect 7472 3612 7524 3664
rect 8484 3612 8536 3664
rect 15200 3612 15252 3664
rect 19064 3612 19116 3664
rect 23388 3612 23440 3664
rect 2228 3408 2280 3460
rect 4804 3544 4856 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5264 3544 5316 3596
rect 4160 3476 4212 3528
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 7012 3476 7064 3528
rect 7656 3476 7708 3528
rect 8024 3476 8076 3528
rect 8484 3476 8536 3528
rect 10876 3544 10928 3596
rect 12072 3544 12124 3596
rect 17684 3544 17736 3596
rect 9588 3476 9640 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 6276 3340 6328 3392
rect 6644 3340 6696 3392
rect 11796 3476 11848 3528
rect 12532 3476 12584 3528
rect 14280 3476 14332 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 20168 3476 20220 3528
rect 10692 3408 10744 3460
rect 12808 3451 12860 3460
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 12808 3408 12860 3417
rect 14004 3408 14056 3460
rect 18788 3408 18840 3460
rect 23296 3476 23348 3528
rect 25044 3476 25096 3528
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 8944 3340 8996 3392
rect 14740 3340 14792 3392
rect 15476 3340 15528 3392
rect 16488 3340 16540 3392
rect 20996 3340 21048 3392
rect 21088 3340 21140 3392
rect 25228 3340 25280 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 4252 3136 4304 3188
rect 4436 3136 4488 3188
rect 6736 3179 6788 3188
rect 6736 3145 6745 3179
rect 6745 3145 6779 3179
rect 6779 3145 6788 3179
rect 6736 3136 6788 3145
rect 10140 3136 10192 3188
rect 15568 3136 15620 3188
rect 17592 3136 17644 3188
rect 2596 3000 2648 3052
rect 3424 3043 3476 3052
rect 3424 3009 3433 3043
rect 3433 3009 3467 3043
rect 3467 3009 3476 3043
rect 3424 3000 3476 3009
rect 3976 3000 4028 3052
rect 5172 3000 5224 3052
rect 5448 3000 5500 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7748 3000 7800 3052
rect 8944 3000 8996 3052
rect 10232 3000 10284 3052
rect 11704 3068 11756 3120
rect 15016 3068 15068 3120
rect 16580 3068 16632 3120
rect 21088 3136 21140 3188
rect 21180 3136 21232 3188
rect 22100 3136 22152 3188
rect 22192 3179 22244 3188
rect 22192 3145 22201 3179
rect 22201 3145 22235 3179
rect 22235 3145 22244 3179
rect 22192 3136 22244 3145
rect 22836 3136 22888 3188
rect 25044 3179 25096 3188
rect 25044 3145 25053 3179
rect 25053 3145 25087 3179
rect 25087 3145 25096 3179
rect 25044 3136 25096 3145
rect 22744 3111 22796 3120
rect 22744 3077 22753 3111
rect 22753 3077 22787 3111
rect 22787 3077 22796 3111
rect 22744 3068 22796 3077
rect 22928 3111 22980 3120
rect 22928 3077 22937 3111
rect 22937 3077 22971 3111
rect 22971 3077 22980 3111
rect 22928 3068 22980 3077
rect 24584 3111 24636 3120
rect 24584 3077 24593 3111
rect 24593 3077 24627 3111
rect 24627 3077 24636 3111
rect 24584 3068 24636 3077
rect 24768 3068 24820 3120
rect 1860 2864 1912 2916
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 17132 3000 17184 3052
rect 19892 3043 19944 3052
rect 19892 3009 19901 3043
rect 19901 3009 19935 3043
rect 19935 3009 19944 3043
rect 19892 3000 19944 3009
rect 22284 3000 22336 3052
rect 23388 3000 23440 3052
rect 11060 2932 11112 2984
rect 11612 2932 11664 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 21364 2932 21416 2984
rect 23572 2932 23624 2984
rect 8760 2864 8812 2916
rect 5448 2796 5500 2848
rect 11980 2796 12032 2848
rect 16028 2864 16080 2916
rect 23480 2864 23532 2916
rect 24124 3000 24176 3052
rect 24492 2864 24544 2916
rect 15936 2796 15988 2848
rect 19892 2796 19944 2848
rect 22376 2796 22428 2848
rect 23388 2796 23440 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 4160 2592 4212 2644
rect 9128 2592 9180 2644
rect 13912 2592 13964 2644
rect 14372 2592 14424 2644
rect 16488 2592 16540 2644
rect 18880 2592 18932 2644
rect 20444 2592 20496 2644
rect 23204 2592 23256 2644
rect 23664 2592 23716 2644
rect 9680 2524 9732 2576
rect 2780 2456 2832 2508
rect 1860 2388 1912 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 5264 2456 5316 2508
rect 5356 2388 5408 2440
rect 8852 2456 8904 2508
rect 12164 2524 12216 2576
rect 8300 2388 8352 2440
rect 10968 2456 11020 2508
rect 15752 2524 15804 2576
rect 16120 2524 16172 2576
rect 22192 2524 22244 2576
rect 2964 2320 3016 2372
rect 7840 2320 7892 2372
rect 7104 2252 7156 2304
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9956 2388 10008 2440
rect 14372 2456 14424 2508
rect 15108 2456 15160 2508
rect 11888 2388 11940 2440
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 14096 2388 14148 2440
rect 16764 2388 16816 2440
rect 16948 2388 17000 2440
rect 20904 2456 20956 2508
rect 19064 2388 19116 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19524 2388 19576 2440
rect 24768 2456 24820 2508
rect 24124 2388 24176 2440
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 12348 2320 12400 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 16304 2320 16356 2372
rect 24584 2295 24636 2304
rect 24584 2261 24593 2295
rect 24593 2261 24627 2295
rect 24627 2261 24636 2295
rect 24584 2252 24636 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 2872 2048 2924 2100
rect 9772 2048 9824 2100
rect 8300 1980 8352 2032
rect 20536 1980 20588 2032
rect 7656 1912 7708 1964
rect 24584 1912 24636 1964
rect 10968 1844 11020 1896
rect 22100 1844 22152 1896
rect 7104 1776 7156 1828
rect 11336 1776 11388 1828
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 12070 56200 12126 57000
rect 12176 56222 12388 56250
rect 1044 53650 1072 56200
rect 2424 54262 2452 56200
rect 2412 54256 2464 54262
rect 2412 54198 2464 54204
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 3804 53650 3832 56200
rect 5184 54262 5212 56200
rect 5172 54256 5224 54262
rect 5172 54198 5224 54204
rect 4988 54188 5040 54194
rect 4988 54130 5040 54136
rect 6000 54188 6052 54194
rect 6000 54130 6052 54136
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3792 53644 3844 53650
rect 3792 53586 3844 53592
rect 5000 53242 5028 54130
rect 5356 53576 5408 53582
rect 5356 53518 5408 53524
rect 4988 53236 5040 53242
rect 4988 53178 5040 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 5368 52698 5396 53518
rect 5540 53508 5592 53514
rect 5540 53450 5592 53456
rect 5356 52692 5408 52698
rect 5356 52634 5408 52640
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 5552 50522 5580 53450
rect 6012 51542 6040 54130
rect 6564 53650 6592 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7852 54126 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8392 54188 8444 54194
rect 8392 54130 8444 54136
rect 7840 54120 7892 54126
rect 7840 54062 7892 54068
rect 6552 53644 6604 53650
rect 6552 53586 6604 53592
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7564 53100 7616 53106
rect 7564 53042 7616 53048
rect 6000 51536 6052 51542
rect 6000 51478 6052 51484
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 6644 50516 6696 50522
rect 6644 50458 6696 50464
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 6656 48890 6684 50458
rect 7576 50454 7604 53042
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 8404 51610 8432 54130
rect 9324 54126 9352 56200
rect 9588 54188 9640 54194
rect 9588 54130 9640 54136
rect 9312 54120 9364 54126
rect 9312 54062 9364 54068
rect 8484 54052 8536 54058
rect 8484 53994 8536 54000
rect 8392 51604 8444 51610
rect 8392 51546 8444 51552
rect 7840 51400 7892 51406
rect 7840 51342 7892 51348
rect 7564 50448 7616 50454
rect 7564 50390 7616 50396
rect 6644 48884 6696 48890
rect 6644 48826 6696 48832
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 7852 46170 7880 51342
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 8496 50522 8524 53994
rect 9220 53576 9272 53582
rect 9220 53518 9272 53524
rect 9232 51610 9260 53518
rect 9404 52488 9456 52494
rect 9404 52430 9456 52436
rect 9220 51604 9272 51610
rect 9220 51546 9272 51552
rect 8484 50516 8536 50522
rect 8484 50458 8536 50464
rect 8496 50318 8524 50458
rect 8484 50312 8536 50318
rect 8484 50254 8536 50260
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 8496 47734 8524 50254
rect 8668 48816 8720 48822
rect 8668 48758 8720 48764
rect 8680 48550 8708 48758
rect 8852 48612 8904 48618
rect 8852 48554 8904 48560
rect 8668 48544 8720 48550
rect 8668 48486 8720 48492
rect 8484 47728 8536 47734
rect 8484 47670 8536 47676
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7840 46164 7892 46170
rect 7840 46106 7892 46112
rect 8576 45960 8628 45966
rect 8576 45902 8628 45908
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8588 38010 8616 45902
rect 8680 44742 8708 48486
rect 8864 47462 8892 48554
rect 9416 47802 9444 52430
rect 9600 50522 9628 54130
rect 10704 53718 10732 56200
rect 12084 56114 12112 56200
rect 12176 56114 12204 56222
rect 12084 56086 12204 56114
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53712 10744 53718
rect 10692 53654 10744 53660
rect 10692 53576 10744 53582
rect 10692 53518 10744 53524
rect 10416 51400 10468 51406
rect 10416 51342 10468 51348
rect 10324 51332 10376 51338
rect 10324 51274 10376 51280
rect 9588 50516 9640 50522
rect 9588 50458 9640 50464
rect 9496 50448 9548 50454
rect 9496 50390 9548 50396
rect 9508 48142 9536 50390
rect 9588 50312 9640 50318
rect 9588 50254 9640 50260
rect 9496 48136 9548 48142
rect 9496 48078 9548 48084
rect 9404 47796 9456 47802
rect 9404 47738 9456 47744
rect 8852 47456 8904 47462
rect 8852 47398 8904 47404
rect 9128 47456 9180 47462
rect 9128 47398 9180 47404
rect 9140 45082 9168 47398
rect 9416 47054 9444 47738
rect 9404 47048 9456 47054
rect 9404 46990 9456 46996
rect 9416 45554 9444 46990
rect 9508 46034 9536 48078
rect 9496 46028 9548 46034
rect 9496 45970 9548 45976
rect 9232 45526 9444 45554
rect 9128 45076 9180 45082
rect 9128 45018 9180 45024
rect 8668 44736 8720 44742
rect 8668 44678 8720 44684
rect 9232 44402 9260 45526
rect 9600 44538 9628 50254
rect 10232 49156 10284 49162
rect 10232 49098 10284 49104
rect 9772 46708 9824 46714
rect 9772 46650 9824 46656
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 8944 44328 8996 44334
rect 8944 44270 8996 44276
rect 8576 38004 8628 38010
rect 8576 37946 8628 37952
rect 8852 37868 8904 37874
rect 8852 37810 8904 37816
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23662 7880 24142
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8404 23798 8432 24006
rect 8392 23792 8444 23798
rect 8392 23734 8444 23740
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6932 21486 6960 22102
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 6932 20466 6960 21422
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 6564 19310 6592 20402
rect 7576 19310 7604 22714
rect 7852 22166 7880 23598
rect 8208 23248 8260 23254
rect 8208 23190 8260 23196
rect 8220 22964 8248 23190
rect 8220 22936 8340 22964
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8312 22778 8340 22936
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8404 22658 8432 23734
rect 8312 22642 8432 22658
rect 8300 22636 8432 22642
rect 8352 22630 8432 22636
rect 8300 22578 8352 22584
rect 7840 22160 7892 22166
rect 7840 22102 7892 22108
rect 8312 21894 8340 22578
rect 8496 22094 8524 26250
rect 8404 22066 8524 22094
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8312 21554 8340 21830
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7760 19258 7788 21422
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20534 8340 21490
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8312 19718 8340 20470
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8208 19440 8260 19446
rect 8312 19428 8340 19654
rect 8260 19400 8340 19428
rect 8208 19382 8260 19388
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 6564 18766 6592 19246
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6564 18426 6592 18702
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 6564 16114 6592 18362
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 6840 15502 6868 15982
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 6564 13530 6592 15438
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14346 6868 14894
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6840 13938 6868 14282
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6932 12918 6960 19246
rect 7760 19242 7880 19258
rect 7760 19236 7892 19242
rect 7760 19230 7840 19236
rect 7760 18222 7788 19230
rect 7840 19178 7892 19184
rect 8220 18714 8248 19382
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18834 8340 19110
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8220 18698 8340 18714
rect 8220 18692 8352 18698
rect 8220 18686 8300 18692
rect 8300 18634 8352 18640
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8208 18352 8260 18358
rect 8312 18340 8340 18634
rect 8260 18312 8340 18340
rect 8208 18294 8260 18300
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17338 7420 17478
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7300 13394 7328 14418
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3896 8809 3924 9590
rect 3882 8800 3938 8809
rect 3882 8735 3938 8744
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1504 3398 1532 4082
rect 1596 3738 1624 4558
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 2688 3936 2740 3942
rect 3424 3936 3476 3942
rect 2740 3896 2820 3924
rect 2688 3878 2740 3884
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 800 1532 3334
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1872 2446 1900 2858
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1872 800 1900 2382
rect 2240 800 2268 3402
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 800 2636 2994
rect 2792 2514 2820 3896
rect 3424 3878 3476 3884
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3436 3058 3464 3878
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3436 2774 3464 2994
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2746 3464 2774
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2884 2106 2912 2382
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2976 800 3004 2314
rect 3344 800 3372 2746
rect 3712 800 3740 3946
rect 3988 3058 4016 11494
rect 5354 9208 5410 9217
rect 5354 9143 5410 9152
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6497 4108 6598
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4080 3942 4108 4082
rect 5170 4040 5226 4049
rect 5170 3975 5226 3984
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4080 800 4108 3878
rect 5184 3602 5212 3975
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3602 5304 3878
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4172 2650 4200 3470
rect 4264 3194 4292 3470
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4448 800 4476 3130
rect 4816 800 4844 3538
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5184 800 5212 2994
rect 5368 2774 5396 9143
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5920 4010 5948 4082
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3058 5488 3878
rect 5722 3088 5778 3097
rect 5448 3052 5500 3058
rect 5722 3023 5778 3032
rect 5448 2994 5500 3000
rect 5736 2990 5764 3023
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5276 2746 5396 2774
rect 5276 2514 5304 2746
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5356 2440 5408 2446
rect 5460 2428 5488 2790
rect 5408 2400 5488 2428
rect 5356 2382 5408 2388
rect 5460 1714 5488 2400
rect 5460 1686 5580 1714
rect 5552 800 5580 1686
rect 5920 800 5948 3946
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 800 6316 3334
rect 6564 3058 6592 3946
rect 6656 3398 6684 6258
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6748 3194 6776 6122
rect 7024 4078 7052 12650
rect 7300 12238 7328 13330
rect 7392 13002 7420 17138
rect 7392 12974 7512 13002
rect 7576 12986 7604 18022
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7668 13530 7696 17546
rect 7852 14618 7880 17682
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16182 8340 18312
rect 8404 17134 8432 22066
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16794 8432 17070
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8312 14958 8340 15846
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 13852 7880 14554
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8024 13864 8076 13870
rect 7852 13824 8024 13852
rect 8024 13806 8076 13812
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 8312 13326 8340 13942
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7392 12306 7420 12786
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7300 11898 7328 12174
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 9722 7144 10406
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7116 4622 7144 9658
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7024 3534 7052 3878
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6564 2774 6592 2994
rect 6564 2746 6684 2774
rect 6656 800 6684 2746
rect 7024 800 7052 3470
rect 7208 3058 7236 3878
rect 7484 3670 7512 12974
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7208 2774 7236 2994
rect 7208 2746 7420 2774
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1834 7144 2246
rect 7104 1828 7156 1834
rect 7104 1770 7156 1776
rect 7392 800 7420 2746
rect 7668 1970 7696 3470
rect 7760 3058 7788 3878
rect 7852 3738 7880 12786
rect 8220 12306 8248 12786
rect 8496 12782 8524 18906
rect 8588 17882 8616 30194
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8680 21690 8708 23122
rect 8668 21684 8720 21690
rect 8668 21626 8720 21632
rect 8680 20398 8708 21626
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8772 19514 8800 30670
rect 8864 29306 8892 37810
rect 8956 34202 8984 44270
rect 9784 42770 9812 46650
rect 10244 42770 10272 49098
rect 10336 46714 10364 51274
rect 10324 46708 10376 46714
rect 10324 46650 10376 46656
rect 10428 45966 10456 51342
rect 10704 49366 10732 53518
rect 11716 49366 11744 54130
rect 12360 54126 12388 56222
rect 13450 56200 13506 57000
rect 13556 56222 13768 56250
rect 13464 56114 13492 56200
rect 13556 56114 13584 56222
rect 13464 56086 13584 56114
rect 13740 55214 13768 56222
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 16316 56222 16528 56250
rect 13740 55186 13860 55214
rect 13832 54330 13860 55186
rect 13820 54324 13872 54330
rect 13820 54266 13872 54272
rect 14844 54194 14872 56200
rect 16224 56114 16252 56200
rect 16316 56114 16344 56222
rect 16224 56086 16344 56114
rect 14832 54188 14884 54194
rect 16500 54176 16528 56222
rect 17590 56200 17646 57000
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 20456 56222 20668 56250
rect 17604 54194 17632 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18984 54330 19012 56200
rect 20364 56114 20392 56200
rect 20456 56114 20484 56222
rect 20364 56086 20484 56114
rect 18972 54324 19024 54330
rect 18972 54266 19024 54272
rect 16580 54188 16632 54194
rect 16500 54148 16580 54176
rect 14832 54130 14884 54136
rect 16580 54130 16632 54136
rect 17592 54188 17644 54194
rect 20640 54176 20668 56222
rect 21730 56200 21786 57000
rect 21836 56222 22048 56250
rect 21744 56114 21772 56200
rect 21836 56114 21864 56222
rect 21744 56086 21864 56114
rect 20720 54188 20772 54194
rect 20640 54148 20720 54176
rect 17592 54130 17644 54136
rect 22020 54176 22048 56222
rect 23110 56200 23166 57000
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 23124 55214 23152 56200
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 23124 55186 23336 55214
rect 22100 54188 22152 54194
rect 22020 54148 22100 54176
rect 20720 54130 20772 54136
rect 22100 54130 22152 54136
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 13912 54052 13964 54058
rect 13912 53994 13964 54000
rect 16764 54052 16816 54058
rect 16764 53994 16816 54000
rect 12716 53984 12768 53990
rect 12716 53926 12768 53932
rect 10692 49360 10744 49366
rect 10692 49302 10744 49308
rect 11704 49360 11756 49366
rect 11704 49302 11756 49308
rect 10968 49156 11020 49162
rect 10968 49098 11020 49104
rect 10876 48544 10928 48550
rect 10876 48486 10928 48492
rect 10784 47728 10836 47734
rect 10784 47670 10836 47676
rect 10796 46714 10824 47670
rect 10784 46708 10836 46714
rect 10784 46650 10836 46656
rect 10796 46578 10824 46650
rect 10784 46572 10836 46578
rect 10784 46514 10836 46520
rect 10600 46368 10652 46374
rect 10600 46310 10652 46316
rect 10416 45960 10468 45966
rect 10416 45902 10468 45908
rect 10428 44198 10456 45902
rect 10612 44810 10640 46310
rect 10888 44878 10916 48486
rect 10876 44872 10928 44878
rect 10876 44814 10928 44820
rect 10600 44804 10652 44810
rect 10600 44746 10652 44752
rect 10416 44192 10468 44198
rect 10416 44134 10468 44140
rect 9772 42764 9824 42770
rect 9772 42706 9824 42712
rect 10232 42764 10284 42770
rect 10232 42706 10284 42712
rect 9036 42696 9088 42702
rect 9036 42638 9088 42644
rect 8944 34196 8996 34202
rect 8944 34138 8996 34144
rect 9048 30122 9076 42638
rect 10428 41682 10456 44134
rect 10612 42362 10640 44746
rect 10980 44282 11008 49098
rect 12624 48000 12676 48006
rect 12624 47942 12676 47948
rect 11060 46708 11112 46714
rect 11060 46650 11112 46656
rect 11072 44402 11100 46650
rect 12636 45558 12664 47942
rect 12624 45552 12676 45558
rect 12624 45494 12676 45500
rect 12728 45490 12756 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13728 46980 13780 46986
rect 13728 46922 13780 46928
rect 13740 46646 13768 46922
rect 13728 46640 13780 46646
rect 13728 46582 13780 46588
rect 13924 46578 13952 53994
rect 13912 46572 13964 46578
rect 13912 46514 13964 46520
rect 15752 46504 15804 46510
rect 15752 46446 15804 46452
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 15108 45824 15160 45830
rect 15108 45766 15160 45772
rect 12716 45484 12768 45490
rect 12716 45426 12768 45432
rect 14556 45416 14608 45422
rect 14556 45358 14608 45364
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 11152 44736 11204 44742
rect 11152 44678 11204 44684
rect 11336 44736 11388 44742
rect 11336 44678 11388 44684
rect 11060 44396 11112 44402
rect 11060 44338 11112 44344
rect 10888 44254 11008 44282
rect 10600 42356 10652 42362
rect 10600 42298 10652 42304
rect 10888 41818 10916 44254
rect 10968 44192 11020 44198
rect 10968 44134 11020 44140
rect 10980 42294 11008 44134
rect 11164 42362 11192 44678
rect 11152 42356 11204 42362
rect 11152 42298 11204 42304
rect 10968 42288 11020 42294
rect 10968 42230 11020 42236
rect 10876 41812 10928 41818
rect 10876 41754 10928 41760
rect 10416 41676 10468 41682
rect 10416 41618 10468 41624
rect 10232 41608 10284 41614
rect 10232 41550 10284 41556
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 9036 30116 9088 30122
rect 9036 30058 9088 30064
rect 8852 29300 8904 29306
rect 8852 29242 8904 29248
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9140 24070 9168 24754
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9232 23322 9260 33934
rect 9692 29102 9720 35566
rect 10244 30938 10272 41550
rect 10980 35630 11008 42230
rect 11348 42158 11376 44678
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 11520 42356 11572 42362
rect 11520 42298 11572 42304
rect 11336 42152 11388 42158
rect 11336 42094 11388 42100
rect 11532 42022 11560 42298
rect 11520 42016 11572 42022
rect 11520 41958 11572 41964
rect 11704 42016 11756 42022
rect 11704 41958 11756 41964
rect 11532 35766 11560 41958
rect 11716 35894 11744 41958
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 11716 35866 11836 35894
rect 11716 35834 11744 35866
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 11532 30326 11560 35702
rect 11808 35494 11836 35866
rect 11796 35488 11848 35494
rect 11796 35430 11848 35436
rect 11808 34066 11836 35430
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 11796 30048 11848 30054
rect 11796 29990 11848 29996
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11060 29572 11112 29578
rect 11060 29514 11112 29520
rect 10232 29232 10284 29238
rect 10232 29174 10284 29180
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9692 28778 9720 29038
rect 9600 28762 9720 28778
rect 9588 28756 9720 28762
rect 9640 28750 9720 28756
rect 9588 28698 9640 28704
rect 9588 28484 9640 28490
rect 9588 28426 9640 28432
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9324 26858 9352 27270
rect 9600 27130 9628 28426
rect 9864 27940 9916 27946
rect 9864 27882 9916 27888
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9876 27062 9904 27882
rect 9864 27056 9916 27062
rect 9864 26998 9916 27004
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9232 20806 9260 21490
rect 9324 21486 9352 26794
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9416 26314 9444 26522
rect 9876 26450 9904 26998
rect 9864 26444 9916 26450
rect 9864 26386 9916 26392
rect 9404 26308 9456 26314
rect 9404 26250 9456 26256
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9692 24834 9720 25094
rect 9508 24806 9720 24834
rect 9404 24608 9456 24614
rect 9404 24550 9456 24556
rect 9416 24410 9444 24550
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9508 24138 9536 24806
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8588 15910 8616 16118
rect 8680 15978 8708 19246
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8588 15178 8616 15846
rect 8588 15150 8708 15178
rect 8680 15094 8708 15150
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8680 14278 8708 15030
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 14006 8708 14214
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8680 13190 8708 13942
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8680 11898 8708 13126
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8036 3534 8064 3878
rect 8496 3670 8524 10542
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8588 3738 8616 7754
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8024 3528 8076 3534
rect 7930 3496 7986 3505
rect 8024 3470 8076 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 7930 3431 7986 3440
rect 7944 3398 7972 3431
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7656 1964 7708 1970
rect 7656 1906 7708 1912
rect 7760 800 7788 2994
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 2314
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8312 2038 8340 2382
rect 8300 2032 8352 2038
rect 8300 1974 8352 1980
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 3470
rect 8772 2922 8800 18566
rect 8864 9654 8892 18634
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8956 12850 8984 17138
rect 9048 15706 9076 19314
rect 9140 18426 9168 19790
rect 9232 18630 9260 20742
rect 9416 19922 9444 22374
rect 9404 19916 9456 19922
rect 9324 19876 9404 19904
rect 9324 18970 9352 19876
rect 9404 19858 9456 19864
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9416 18698 9444 19246
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9508 18442 9536 24074
rect 9600 22710 9628 24346
rect 9588 22704 9640 22710
rect 9588 22646 9640 22652
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9692 22166 9720 22646
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9692 21010 9720 22102
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19514 9628 19654
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9232 18414 9536 18442
rect 9232 17134 9260 18414
rect 9600 18290 9628 19110
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9508 17746 9536 18226
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 17882 9720 18158
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 17338 9444 17478
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9508 17270 9536 17682
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9048 13326 9076 13806
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8956 12102 8984 12786
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8956 4146 8984 12038
rect 9048 11676 9076 13262
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9140 12782 9168 13194
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9128 11688 9180 11694
rect 9048 11648 9128 11676
rect 9128 11630 9180 11636
rect 9140 11150 9168 11630
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10470 9168 11086
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9324 9994 9352 14894
rect 9416 12714 9444 15302
rect 9508 12986 9536 15438
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 13938 9628 14350
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9692 11898 9720 13126
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9600 11778 9628 11834
rect 9600 11750 9720 11778
rect 9692 11558 9720 11750
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10130 9628 10406
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9324 7342 9352 8774
rect 9600 7478 9628 10066
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6254 9352 7278
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9600 5710 9628 7414
rect 9784 6662 9812 22170
rect 9968 21690 9996 25842
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9968 20942 9996 21490
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9876 14226 9904 16390
rect 9968 15162 9996 19314
rect 10060 18902 10088 22918
rect 10244 21690 10272 29174
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10428 23866 10456 29106
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10520 23662 10548 24890
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10520 23322 10548 23598
rect 10796 23526 10824 25094
rect 10980 23662 11008 28426
rect 11072 27130 11100 29514
rect 11336 28960 11388 28966
rect 11336 28902 11388 28908
rect 11348 28490 11376 28902
rect 11440 28558 11468 29650
rect 11520 29096 11572 29102
rect 11520 29038 11572 29044
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11336 28484 11388 28490
rect 11336 28426 11388 28432
rect 11244 27396 11296 27402
rect 11244 27338 11296 27344
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11072 25838 11100 27066
rect 11256 27062 11284 27338
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11256 26790 11284 26998
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11256 26314 11284 26726
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 11256 25294 11284 26250
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11072 24154 11100 24550
rect 11164 24274 11192 24686
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11072 24126 11192 24154
rect 11256 24138 11284 25230
rect 11164 24070 11192 24126
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10416 23044 10468 23050
rect 10416 22986 10468 22992
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10428 20602 10456 22986
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 10152 17746 10180 20334
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18426 10364 18566
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 9876 14198 9996 14226
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 12918 9904 14010
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 10742 9904 11494
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 4690 9628 5646
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9232 4146 9260 4422
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3058 8984 3334
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 8864 800 8892 2450
rect 9140 2446 9168 2586
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9232 800 9260 4082
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 800 9628 3470
rect 9692 2582 9720 4490
rect 9968 2774 9996 14198
rect 10152 13870 10180 14282
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10060 10810 10088 12718
rect 10244 12442 10272 17478
rect 10428 16522 10456 20334
rect 10520 18834 10548 23258
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10520 18698 10548 18770
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 10612 16454 10640 21830
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10796 19242 10824 20266
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10796 18766 10824 19178
rect 10888 18970 10916 23598
rect 10980 21486 11008 23598
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11072 22166 11100 23258
rect 11164 22166 11192 24006
rect 11348 23322 11376 28426
rect 11440 27538 11468 28494
rect 11428 27532 11480 27538
rect 11428 27474 11480 27480
rect 11532 26518 11560 29038
rect 11808 28966 11836 29990
rect 11900 29578 11928 30262
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 12544 29306 12572 31894
rect 12636 29306 12664 32710
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 14464 31408 14516 31414
rect 14464 31350 14516 31356
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13452 31136 13504 31142
rect 13452 31078 13504 31084
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12808 30184 12860 30190
rect 12808 30126 12860 30132
rect 12820 29850 12848 30126
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13464 29850 13492 31078
rect 13556 30258 13584 31214
rect 14476 31142 14504 31350
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 13544 30252 13596 30258
rect 13544 30194 13596 30200
rect 14568 30190 14596 45358
rect 15120 44810 15148 45766
rect 15108 44804 15160 44810
rect 15108 44746 15160 44752
rect 15764 35698 15792 46446
rect 16488 46368 16540 46374
rect 16488 46310 16540 46316
rect 16500 45898 16528 46310
rect 16488 45892 16540 45898
rect 16488 45834 16540 45840
rect 16580 43648 16632 43654
rect 16580 43590 16632 43596
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 16304 33924 16356 33930
rect 16304 33866 16356 33872
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15488 31822 15516 32302
rect 16224 31890 16252 32914
rect 16316 32502 16344 33866
rect 16592 32978 16620 43590
rect 16776 33114 16804 53994
rect 16856 53984 16908 53990
rect 16856 53926 16908 53932
rect 17500 53984 17552 53990
rect 17500 53926 17552 53932
rect 22100 53984 22152 53990
rect 22100 53926 22152 53932
rect 16868 46034 16896 53926
rect 17408 52556 17460 52562
rect 17408 52498 17460 52504
rect 16856 46028 16908 46034
rect 16856 45970 16908 45976
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 16580 32972 16632 32978
rect 16580 32914 16632 32920
rect 16776 32910 16804 33050
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16304 32496 16356 32502
rect 16304 32438 16356 32444
rect 16212 31884 16264 31890
rect 16212 31826 16264 31832
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15488 31278 15516 31758
rect 16224 31482 16252 31826
rect 16212 31476 16264 31482
rect 16212 31418 16264 31424
rect 15476 31272 15528 31278
rect 15476 31214 15528 31220
rect 16316 30938 16344 32438
rect 16684 31686 16712 32506
rect 17040 32224 17092 32230
rect 17040 32166 17092 32172
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16672 31680 16724 31686
rect 16672 31622 16724 31628
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 14832 30660 14884 30666
rect 14832 30602 14884 30608
rect 13636 30184 13688 30190
rect 13636 30126 13688 30132
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 12808 29844 12860 29850
rect 12808 29786 12860 29792
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 13452 29844 13504 29850
rect 13452 29786 13504 29792
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 11796 28960 11848 28966
rect 11796 28902 11848 28908
rect 11520 26512 11572 26518
rect 11520 26454 11572 26460
rect 11612 26512 11664 26518
rect 11612 26454 11664 26460
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10980 20058 11008 20810
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 10980 18834 11008 19994
rect 11164 18850 11192 21898
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11072 18822 11192 18850
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 11072 17338 11100 18822
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 11626 10272 11834
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10428 11218 10456 13126
rect 10520 12442 10548 14962
rect 10704 14958 10732 15506
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10796 12458 10824 12650
rect 10508 12436 10560 12442
rect 10796 12430 10916 12458
rect 10508 12378 10560 12384
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10428 10742 10456 11018
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10428 10470 10456 10678
rect 10612 10538 10640 11222
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10152 3194 10180 10066
rect 10612 9042 10640 10474
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10704 8906 10732 9454
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10230 6216 10286 6225
rect 10230 6151 10286 6160
rect 10244 4146 10272 6151
rect 10336 4690 10364 8026
rect 10704 6798 10732 8842
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 5098 10732 6734
rect 10796 5778 10824 7142
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4690 10640 4966
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10888 3602 10916 12430
rect 10980 12306 11008 12718
rect 11164 12646 11192 18634
rect 11256 18358 11284 22918
rect 11348 20602 11376 22986
rect 11440 21894 11468 25910
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11532 19922 11560 24074
rect 11624 23118 11652 26454
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11716 23186 11744 25434
rect 11796 24880 11848 24886
rect 11796 24822 11848 24828
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11440 19242 11468 19654
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11256 17882 11284 18158
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11256 16726 11284 17818
rect 11348 17610 11376 18226
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11256 14482 11284 16662
rect 11348 16182 11376 17274
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11348 15162 11376 16118
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13258 11284 14214
rect 11348 14006 11376 15098
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11440 13682 11468 19178
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11532 17678 11560 18566
rect 11624 18442 11652 21490
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 19514 11744 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11624 18414 11744 18442
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11624 17338 11652 18226
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11348 13654 11468 13682
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11256 12918 11284 13194
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 11348 11898 11376 13654
rect 11532 13512 11560 17002
rect 11716 15706 11744 18414
rect 11808 16998 11836 24822
rect 11992 24818 12020 28970
rect 12728 28490 12756 29446
rect 13004 29102 13032 29786
rect 13648 29714 13676 30126
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 12992 29096 13044 29102
rect 12992 29038 13044 29044
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12716 28484 12768 28490
rect 12716 28426 12768 28432
rect 12728 28218 12756 28426
rect 13372 28422 13400 28902
rect 13556 28422 13584 29242
rect 13648 29238 13676 29650
rect 13636 29232 13688 29238
rect 13636 29174 13688 29180
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 12084 26586 12112 27950
rect 12728 27606 12756 28154
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12348 27600 12400 27606
rect 12348 27542 12400 27548
rect 12716 27600 12768 27606
rect 12716 27542 12768 27548
rect 12360 26790 12388 27542
rect 12728 27470 12756 27542
rect 12716 27464 12768 27470
rect 12716 27406 12768 27412
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 12084 24750 12112 26522
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11900 18222 11928 23258
rect 12360 22642 12388 24210
rect 12544 24138 12572 26726
rect 12636 26042 12664 27270
rect 12728 27062 12756 27406
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12728 24886 12756 26998
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13372 25838 13400 28358
rect 13556 28218 13584 28358
rect 13544 28212 13596 28218
rect 13544 28154 13596 28160
rect 13452 28008 13504 28014
rect 13452 27950 13504 27956
rect 13464 27878 13492 27950
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 13464 27674 13492 27814
rect 13452 27668 13504 27674
rect 13452 27610 13504 27616
rect 13832 27470 13860 28358
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13924 27402 13952 27814
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12728 24274 12756 24822
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12728 24138 12756 24210
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12360 22114 12388 22578
rect 12544 22166 12572 23462
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12532 22160 12584 22166
rect 12360 22086 12480 22114
rect 12532 22102 12584 22108
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12084 18358 12112 20878
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11440 13484 11560 13512
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11072 11150 11100 11630
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 9994 11008 10406
rect 11072 10266 11100 11086
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11440 7970 11468 13484
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11532 9518 11560 13330
rect 11624 10266 11652 14962
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11716 12986 11744 13806
rect 11808 13258 11836 16390
rect 11900 16250 11928 17614
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 17338 12020 17546
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 12084 17066 12112 17478
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 12176 16250 12204 21558
rect 12452 20466 12480 22086
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12452 19922 12480 20402
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 11900 15978 11928 16186
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11900 15570 11928 15914
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11888 13932 11940 13938
rect 11992 13920 12020 15574
rect 12268 15502 12296 17274
rect 12452 16810 12480 19450
rect 12544 17746 12572 20742
rect 12636 18834 12664 22918
rect 12728 22710 12756 24074
rect 12820 22778 12848 25230
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 12912 24750 12940 25094
rect 13004 24886 13032 25094
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 13464 24750 13492 26318
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13556 23882 13584 27270
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13464 23854 13584 23882
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12728 21690 12756 22646
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20330 12756 21286
rect 12820 20874 12848 22714
rect 13004 22438 13032 23122
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12728 17134 12756 20266
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 20058 13400 23802
rect 13464 23662 13492 23854
rect 13648 23798 13676 26522
rect 14660 25906 14688 28970
rect 14844 28558 14872 30602
rect 15304 30326 15332 30670
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15580 29782 15608 30126
rect 16304 30116 16356 30122
rect 16304 30058 16356 30064
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15568 29776 15620 29782
rect 15568 29718 15620 29724
rect 15844 29708 15896 29714
rect 15844 29650 15896 29656
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15108 29300 15160 29306
rect 15108 29242 15160 29248
rect 14832 28552 14884 28558
rect 14832 28494 14884 28500
rect 14844 27946 14872 28494
rect 14832 27940 14884 27946
rect 14832 27882 14884 27888
rect 14844 26994 14872 27882
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13740 24410 13768 24686
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13740 23798 13768 24346
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13728 23792 13780 23798
rect 13728 23734 13780 23740
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13452 23656 13504 23662
rect 13452 23598 13504 23604
rect 13556 23610 13584 23666
rect 13832 23610 13860 25638
rect 14648 25424 14700 25430
rect 14648 25366 14700 25372
rect 14660 25158 14688 25366
rect 14752 25362 14780 26386
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14752 24342 14780 25298
rect 14844 25226 14872 26930
rect 14936 26246 14964 27406
rect 15120 27062 15148 29242
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14844 24818 14872 25162
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14936 23882 14964 26182
rect 13556 23582 13860 23610
rect 14844 23854 14964 23882
rect 15028 23866 15056 26726
rect 15212 25430 15240 29582
rect 15752 29028 15804 29034
rect 15752 28970 15804 28976
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15396 28014 15424 28562
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 15488 26450 15516 28562
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15580 27334 15608 28358
rect 15568 27328 15620 27334
rect 15566 27296 15568 27305
rect 15620 27296 15622 27305
rect 15566 27231 15622 27240
rect 15764 27062 15792 28970
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15384 25832 15436 25838
rect 15384 25774 15436 25780
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 15212 24818 15240 25366
rect 15396 25242 15424 25774
rect 15304 25214 15424 25242
rect 15304 25158 15332 25214
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15304 24954 15332 25094
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 24721 15240 24754
rect 15198 24712 15254 24721
rect 15198 24647 15254 24656
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 15016 23860 15068 23866
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13556 21350 13584 23462
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22778 14504 22918
rect 14844 22778 14872 23854
rect 15016 23802 15068 23808
rect 14924 23792 14976 23798
rect 14924 23734 14976 23740
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13924 21894 13952 22578
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22098 14136 22374
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12452 16782 12572 16810
rect 12544 16658 12572 16782
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15706 12664 15982
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11940 13892 12020 13920
rect 11888 13874 11940 13880
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 11014 11836 12582
rect 11900 11694 11928 13874
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11992 11898 12020 12378
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 10606 11836 10950
rect 11900 10742 11928 11630
rect 11992 11558 12020 11834
rect 12084 11665 12112 15302
rect 12268 15162 12296 15438
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12268 14634 12296 15098
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12176 14606 12296 14634
rect 12176 14346 12204 14606
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12268 14006 12296 14418
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12176 12594 12204 13194
rect 12268 12986 12296 13942
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12268 12782 12296 12922
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12176 12566 12296 12594
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12070 11656 12126 11665
rect 12070 11591 12126 11600
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11900 10062 11928 10542
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11624 9654 11652 9930
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11520 9376 11572 9382
rect 11624 9330 11652 9590
rect 11572 9324 11652 9330
rect 11520 9318 11652 9324
rect 11532 9302 11652 9318
rect 11532 8838 11560 9302
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11256 7942 11468 7970
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11072 6254 11100 6666
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10980 4690 11008 5170
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11072 3942 11100 5714
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 5137 11192 5170
rect 11150 5128 11206 5137
rect 11150 5063 11206 5072
rect 11150 4584 11206 4593
rect 11150 4519 11206 4528
rect 11164 4282 11192 4519
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11256 4049 11284 7942
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11242 4040 11298 4049
rect 11242 3975 11298 3984
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 9784 2746 9996 2774
rect 10244 2774 10272 2994
rect 10244 2746 10364 2774
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9784 2106 9812 2746
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9968 800 9996 2382
rect 10336 800 10364 2746
rect 10704 800 10732 3402
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10980 1902 11008 2450
rect 10968 1896 11020 1902
rect 10968 1838 11020 1844
rect 11072 800 11100 2926
rect 11348 1834 11376 7686
rect 11532 7478 11560 8774
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11716 7886 11744 8366
rect 11796 8016 11848 8022
rect 11794 7984 11796 7993
rect 11848 7984 11850 7993
rect 11794 7919 11850 7928
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11900 7546 11928 7890
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11532 7274 11560 7414
rect 11900 7274 11928 7482
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6390 11468 7142
rect 11532 6730 11560 7210
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11440 5846 11468 6326
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11428 5704 11480 5710
rect 11532 5658 11560 6666
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5914 11836 6190
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11480 5652 11560 5658
rect 11428 5646 11560 5652
rect 11440 5630 11560 5646
rect 11440 4758 11468 5630
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11624 2990 11652 4422
rect 11808 3534 11836 5238
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11624 2774 11652 2926
rect 11440 2746 11652 2774
rect 11336 1828 11388 1834
rect 11336 1770 11388 1776
rect 11440 800 11468 2746
rect 11716 1442 11744 3062
rect 11900 2446 11928 3878
rect 11992 2854 12020 11494
rect 12176 10130 12204 12242
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12268 7562 12296 12566
rect 12360 10130 12388 13126
rect 12452 12481 12480 14894
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 13938 12572 14758
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12438 12472 12494 12481
rect 12438 12407 12494 12416
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12360 9178 12388 9658
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 9110 12480 12310
rect 12544 12306 12572 12650
rect 12636 12442 12664 15370
rect 12820 14618 12848 18566
rect 13280 18170 13308 18566
rect 13372 18358 13400 19858
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13924 19174 13952 19382
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13360 18352 13412 18358
rect 13412 18312 13584 18340
rect 13360 18294 13412 18300
rect 13452 18216 13504 18222
rect 13280 18142 13400 18170
rect 13452 18158 13504 18164
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17338 13216 17478
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13188 15910 13216 16594
rect 13280 16250 13308 16730
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 12646 12756 13806
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12714 12472 12770 12481
rect 12624 12436 12676 12442
rect 12714 12407 12770 12416
rect 12624 12378 12676 12384
rect 12728 12374 12756 12407
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12544 11082 12572 12106
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11354 12756 12038
rect 12820 11898 12848 14214
rect 13004 14074 13032 14418
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13280 12850 13308 13398
rect 13372 12986 13400 18142
rect 13464 17814 13492 18158
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13464 16538 13492 17750
rect 13556 16658 13584 18312
rect 14016 17882 14044 21830
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14292 19922 14320 21558
rect 14568 21486 14596 22034
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14660 20534 14688 20742
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14292 19378 14320 19858
rect 14476 19446 14504 20198
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14200 18426 14228 18566
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13464 16510 13584 16538
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15638 13492 15914
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13280 12730 13308 12786
rect 13280 12702 13400 12730
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13096 11898 13124 12242
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 13082 11656 13138 11665
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12636 10810 12664 11222
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12728 10810 12756 11018
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12820 10010 12848 11630
rect 13082 11591 13084 11600
rect 13136 11591 13138 11600
rect 13084 11562 13136 11568
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12912 10606 12940 11290
rect 13004 11014 13032 11290
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12544 9982 12848 10010
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12268 7534 12388 7562
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 3602 12112 7346
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 12176 2582 12204 6258
rect 12254 5808 12310 5817
rect 12254 5743 12310 5752
rect 12268 5710 12296 5743
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12254 5400 12310 5409
rect 12254 5335 12310 5344
rect 12268 5234 12296 5335
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11716 1414 11836 1442
rect 11808 800 11836 1414
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 11900 762 11928 2382
rect 12360 2378 12388 7534
rect 12544 7426 12572 9982
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12636 8974 12664 9114
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12728 8022 12756 9454
rect 12820 9178 12848 9862
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13372 8634 13400 12702
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 9926 13492 12582
rect 13556 12442 13584 16510
rect 13648 16046 13676 17070
rect 13832 16182 13860 17750
rect 14200 17610 14228 18362
rect 14292 17678 14320 18566
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14476 16794 14504 19110
rect 14568 18970 14596 19858
rect 14936 19802 14964 23734
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15120 21350 15148 21626
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15120 20534 15148 21286
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15120 20058 15148 20470
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 14844 19786 14964 19802
rect 15120 19786 15148 19994
rect 14832 19780 14964 19786
rect 14884 19774 14964 19780
rect 15108 19780 15160 19786
rect 14832 19722 14884 19728
rect 15108 19722 15160 19728
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 16250 14228 16390
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 13820 16176 13872 16182
rect 13872 16136 13952 16164
rect 13820 16118 13872 16124
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13648 15348 13676 15982
rect 13728 15360 13780 15366
rect 13648 15320 13728 15348
rect 13728 15302 13780 15308
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13648 12322 13676 12786
rect 13556 12294 13676 12322
rect 13556 11898 13584 12294
rect 13740 12186 13768 15302
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 14278 13860 14350
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 13977 13860 14214
rect 13818 13968 13874 13977
rect 13818 13903 13874 13912
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13394 13860 13806
rect 13924 13530 13952 16136
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13924 13326 13952 13466
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 14016 12866 14044 16050
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 13924 12838 14044 12866
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13648 12158 13768 12186
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10130 13584 11154
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 12806 8528 12862 8537
rect 12806 8463 12862 8472
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12452 7398 12572 7426
rect 12452 5778 12480 7398
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12544 6186 12572 7278
rect 12728 6866 12756 7958
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12820 6458 12848 8463
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13372 7886 13400 8366
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 13004 5574 13032 5782
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12898 5264 12954 5273
rect 12898 5199 12900 5208
rect 12952 5199 12954 5208
rect 12900 5170 12952 5176
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12440 4072 12492 4078
rect 12808 4072 12860 4078
rect 12440 4014 12492 4020
rect 12806 4040 12808 4049
rect 12860 4040 12862 4049
rect 12452 2446 12480 4014
rect 12806 3975 12862 3984
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12084 870 12204 898
rect 12084 762 12112 870
rect 12176 800 12204 870
rect 12544 800 12572 3470
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12820 1714 12848 3402
rect 13372 3097 13400 6870
rect 13464 5710 13492 9862
rect 13556 9042 13584 10066
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13542 8936 13598 8945
rect 13542 8871 13544 8880
rect 13596 8871 13598 8880
rect 13544 8842 13596 8848
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13556 6254 13584 7142
rect 13648 6934 13676 12158
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10266 13768 10542
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9450 13768 9930
rect 13832 9518 13860 12718
rect 13924 12594 13952 12838
rect 14004 12776 14056 12782
rect 14108 12764 14136 13670
rect 14056 12736 14136 12764
rect 14004 12718 14056 12724
rect 13924 12566 14136 12594
rect 14108 12442 14136 12566
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11286 13952 12038
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13832 7410 13860 8842
rect 13924 8430 13952 10542
rect 14016 9518 14044 12242
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14108 10441 14136 11154
rect 14200 10810 14228 14282
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14278 12472 14334 12481
rect 14278 12407 14334 12416
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14094 10432 14150 10441
rect 14094 10367 14150 10376
rect 14200 10198 14228 10610
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13728 6792 13780 6798
rect 13634 6760 13690 6769
rect 13728 6734 13780 6740
rect 13634 6695 13690 6704
rect 13648 6662 13676 6695
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13556 5302 13584 6190
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13740 4622 13768 6734
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13832 5914 13860 6326
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13924 5794 13952 8366
rect 13832 5766 13952 5794
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13358 3088 13414 3097
rect 13358 3023 13414 3032
rect 13464 2961 13492 4082
rect 13832 3738 13860 5766
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13924 4146 13952 4966
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14016 4026 14044 9046
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14108 8090 14136 8570
rect 14200 8090 14228 8774
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14094 6488 14150 6497
rect 14094 6423 14150 6432
rect 14108 6254 14136 6423
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 13924 3998 14044 4026
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13636 2984 13688 2990
rect 13450 2952 13506 2961
rect 13636 2926 13688 2932
rect 13450 2887 13506 2896
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 1686 12940 1714
rect 12912 800 12940 1686
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 13924 2650 13952 3998
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14016 800 14044 3402
rect 14108 2446 14136 5782
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4214 14228 4966
rect 14292 4826 14320 12407
rect 14384 11830 14412 14214
rect 14476 11898 14504 15642
rect 14568 14958 14596 17070
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14568 12986 14596 13466
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14476 11082 14504 11222
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14476 9518 14504 10066
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14384 9382 14412 9454
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8498 14412 9318
rect 14476 9042 14504 9454
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8566 14504 8978
rect 14568 8838 14596 11698
rect 14660 11558 14688 19178
rect 14844 17134 14872 19722
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15028 18154 15056 19314
rect 15120 19174 15148 19722
rect 15212 19514 15240 20946
rect 15396 20602 15424 24618
rect 15488 24614 15516 26386
rect 15856 25226 15884 29650
rect 15948 29306 15976 29990
rect 16316 29850 16344 30058
rect 16304 29844 16356 29850
rect 16304 29786 16356 29792
rect 16316 29646 16344 29786
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16592 29578 16620 31078
rect 16580 29572 16632 29578
rect 16580 29514 16632 29520
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16040 29306 16068 29446
rect 15936 29300 15988 29306
rect 15936 29242 15988 29248
rect 16028 29300 16080 29306
rect 16028 29242 16080 29248
rect 16592 29050 16620 29514
rect 16408 29022 16620 29050
rect 16408 28626 16436 29022
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16408 28490 16436 28562
rect 16396 28484 16448 28490
rect 16396 28426 16448 28432
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 16304 28416 16356 28422
rect 16304 28358 16356 28364
rect 16132 28121 16160 28358
rect 16118 28112 16174 28121
rect 16118 28047 16174 28056
rect 16132 27334 16160 28047
rect 16212 27532 16264 27538
rect 16212 27474 16264 27480
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15844 25220 15896 25226
rect 15844 25162 15896 25168
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15488 24274 15516 24550
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15672 23118 15700 23598
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15764 22166 15792 25094
rect 15856 24818 15884 25162
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15948 22234 15976 26998
rect 16224 26450 16252 27474
rect 16316 27334 16344 28358
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16212 26444 16264 26450
rect 16212 26386 16264 26392
rect 16316 25158 16344 27270
rect 16408 26586 16436 28154
rect 16500 28082 16528 28902
rect 16684 28150 16712 31622
rect 16776 31346 16804 31758
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16868 31142 16896 31962
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16672 28144 16724 28150
rect 16672 28086 16724 28092
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16500 27418 16528 28018
rect 16672 27940 16724 27946
rect 16672 27882 16724 27888
rect 16500 27390 16620 27418
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16396 26580 16448 26586
rect 16396 26522 16448 26528
rect 16408 26314 16436 26522
rect 16396 26308 16448 26314
rect 16396 26250 16448 26256
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16500 24698 16528 27270
rect 16592 26518 16620 27390
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16408 24670 16528 24698
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15856 21554 15884 21830
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15948 21434 15976 21898
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15856 21406 15976 21434
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 15396 17338 15424 20402
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14844 16250 14872 16390
rect 14936 16250 14964 16390
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15366 14780 16050
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15638 15056 15982
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14752 14414 14780 15302
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15212 14482 15240 14962
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15200 14476 15252 14482
rect 15252 14436 15332 14464
rect 15200 14418 15252 14424
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14752 12481 14780 14010
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 15212 13274 15240 13738
rect 15304 13394 15332 14436
rect 15396 14346 15424 14486
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14936 13190 14964 13262
rect 15212 13246 15332 13274
rect 15488 13258 15516 14758
rect 15580 13462 15608 21354
rect 15856 20806 15884 21406
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 19446 15792 20198
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 16590 15700 17478
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15764 16794 15792 17274
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15856 16658 15884 20742
rect 16408 19378 16436 24670
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16500 21962 16528 24550
rect 16684 24070 16712 27882
rect 16776 27470 16804 30126
rect 16960 30054 16988 30194
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16960 29850 16988 29990
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16776 26450 16804 27406
rect 16868 27130 16896 27814
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16960 26450 16988 29786
rect 17052 27946 17080 32166
rect 17132 31748 17184 31754
rect 17132 31690 17184 31696
rect 17144 31482 17172 31690
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 17144 30938 17172 31418
rect 17132 30932 17184 30938
rect 17132 30874 17184 30880
rect 17236 29170 17264 32710
rect 17328 31754 17356 33050
rect 17420 32026 17448 52498
rect 17512 44946 17540 53926
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 21824 48000 21876 48006
rect 21824 47942 21876 47948
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 21732 46096 21784 46102
rect 21732 46038 21784 46044
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 19984 45008 20036 45014
rect 19984 44950 20036 44956
rect 17500 44940 17552 44946
rect 17500 44882 17552 44888
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 19248 35556 19300 35562
rect 19248 35498 19300 35504
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17776 31884 17828 31890
rect 17776 31826 17828 31832
rect 17328 31726 17448 31754
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17328 28082 17356 31078
rect 17420 29306 17448 31726
rect 17788 31278 17816 31826
rect 18788 31680 18840 31686
rect 18788 31622 18840 31628
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18800 31346 18828 31622
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 17776 31272 17828 31278
rect 17776 31214 17828 31220
rect 17684 31136 17736 31142
rect 17684 31078 17736 31084
rect 17696 30818 17724 31078
rect 17604 30790 17724 30818
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17420 29186 17448 29242
rect 17420 29158 17540 29186
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17316 28076 17368 28082
rect 17316 28018 17368 28024
rect 17420 28014 17448 29038
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17040 27940 17092 27946
rect 17040 27882 17092 27888
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 17132 26512 17184 26518
rect 17132 26454 17184 26460
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16776 24070 16804 26386
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16868 25906 16896 25978
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 17052 25362 17080 25638
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16960 24750 16988 25230
rect 17144 24834 17172 26454
rect 17236 24954 17264 26522
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17144 24806 17264 24834
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16592 20058 16620 20810
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15948 15450 15976 17206
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15856 15422 15976 15450
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13530 15700 14214
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14738 12472 14794 12481
rect 14844 12442 14872 12922
rect 14738 12407 14794 12416
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14752 11898 14780 12242
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11694 14872 12242
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14648 11552 14700 11558
rect 14646 11520 14648 11529
rect 14700 11520 14702 11529
rect 14646 11455 14702 11464
rect 14752 10062 14780 11630
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14752 9058 14780 9998
rect 14844 9450 14872 11086
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14752 9030 14872 9058
rect 14844 8906 14872 9030
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14372 8492 14424 8498
rect 14936 8480 14964 13126
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 8650 15056 10950
rect 15120 10130 15148 12310
rect 15212 11354 15240 13126
rect 15304 12866 15332 13246
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15488 12986 15516 13194
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15568 12912 15620 12918
rect 15304 12838 15516 12866
rect 15568 12854 15620 12860
rect 15488 12782 15516 12838
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15304 12442 15332 12718
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15396 12617 15424 12650
rect 15382 12608 15438 12617
rect 15382 12543 15438 12552
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15488 12374 15516 12718
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 11234 15332 11494
rect 15212 11206 15332 11234
rect 15212 11082 15240 11206
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15028 8622 15148 8650
rect 14372 8434 14424 8440
rect 14752 8452 14964 8480
rect 15016 8492 15068 8498
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14370 6896 14426 6905
rect 14476 6866 14504 7414
rect 14370 6831 14426 6840
rect 14464 6860 14516 6866
rect 14384 6662 14412 6831
rect 14464 6802 14516 6808
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14476 6118 14504 6802
rect 14568 6186 14596 7686
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 6186 14688 6666
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5642 14504 6054
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14476 5302 14504 5578
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14292 3534 14320 4762
rect 14370 4040 14426 4049
rect 14370 3975 14426 3984
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14384 3058 14412 3975
rect 14752 3398 14780 8452
rect 15016 8434 15068 8440
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14844 3058 14872 8298
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14936 4690 14964 5102
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 15028 3126 15056 8434
rect 15120 7342 15148 8622
rect 15212 7954 15240 11018
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10470 15332 10542
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 9722 15332 10406
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15396 9586 15424 12038
rect 15580 10810 15608 12854
rect 15764 12764 15792 13466
rect 15672 12736 15792 12764
rect 15672 11898 15700 12736
rect 15750 12608 15806 12617
rect 15750 12543 15806 12552
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15488 10674 15516 10746
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15580 10010 15608 10202
rect 15488 9982 15608 10010
rect 15488 9926 15516 9982
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 8838 15424 9522
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15304 7750 15332 8774
rect 15396 8362 15424 8774
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15488 7562 15516 9658
rect 15580 8838 15608 9862
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15672 9110 15700 9454
rect 15764 9178 15792 12543
rect 15856 12102 15884 15422
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15948 15162 15976 15302
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 16040 14482 16068 17070
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 15910 16160 16390
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16040 14074 16068 14418
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15948 11370 15976 13330
rect 16132 13326 16160 15846
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 15856 11342 15976 11370
rect 15856 9518 15884 11342
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15212 7534 15516 7562
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15212 3670 15240 7534
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15290 5672 15346 5681
rect 15290 5607 15346 5616
rect 15304 5574 15332 5607
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15304 4554 15332 5238
rect 15396 4554 15424 5714
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15396 4298 15424 4490
rect 15396 4282 15516 4298
rect 15396 4276 15528 4282
rect 15396 4270 15476 4276
rect 15476 4218 15528 4224
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14384 2650 14412 2994
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14384 800 14412 2450
rect 14752 800 14780 2926
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15120 800 15148 2450
rect 15488 800 15516 3334
rect 15580 3194 15608 8774
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 4010 15700 8366
rect 15856 7954 15884 9454
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 5166 15884 7686
rect 15948 7342 15976 11154
rect 16040 10606 16068 12310
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16040 9926 16068 10202
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16132 9654 16160 10542
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16040 8974 16068 9454
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15948 6866 15976 7278
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 5710 15976 6802
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15658 3632 15714 3641
rect 15658 3567 15714 3576
rect 15672 3534 15700 3567
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15764 2582 15792 5102
rect 15948 4690 15976 5646
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16040 4570 16068 8910
rect 16120 8424 16172 8430
rect 16224 8401 16252 16934
rect 16316 15162 16344 17546
rect 16408 15706 16436 18770
rect 16500 16454 16528 19654
rect 16592 19310 16620 19994
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16592 16130 16620 18362
rect 16684 17814 16712 24006
rect 16776 23866 16804 24006
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 17052 23730 17080 24686
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16960 21010 16988 22034
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16776 20262 16804 20538
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 18222 16804 20198
rect 16856 18284 16908 18290
rect 16960 18272 16988 20946
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 20058 17080 20198
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17144 19514 17172 23462
rect 17236 20942 17264 24806
rect 17328 23526 17356 26250
rect 17408 25832 17460 25838
rect 17406 25800 17408 25809
rect 17460 25800 17462 25809
rect 17406 25735 17462 25744
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17316 23316 17368 23322
rect 17316 23258 17368 23264
rect 17328 22817 17356 23258
rect 17314 22808 17370 22817
rect 17314 22743 17370 22752
rect 17420 22094 17448 25638
rect 17512 23866 17540 29158
rect 17604 27334 17632 30790
rect 17684 29028 17736 29034
rect 17684 28970 17736 28976
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17604 25294 17632 25706
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17328 22066 17448 22094
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17236 20466 17264 20742
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17236 19990 17264 20402
rect 17224 19984 17276 19990
rect 17224 19926 17276 19932
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16908 18244 16988 18272
rect 16856 18226 16908 18232
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16684 16522 16712 17750
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16684 16250 16712 16458
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16592 16102 16712 16130
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16408 11558 16436 15642
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16500 11830 16528 13806
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16316 10810 16344 11290
rect 16500 11286 16528 11630
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16316 9042 16344 9590
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16120 8366 16172 8372
rect 16210 8392 16266 8401
rect 16132 7886 16160 8366
rect 16210 8327 16266 8336
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16224 7750 16252 8230
rect 16408 7818 16436 9862
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16316 6934 16344 7754
rect 16500 7478 16528 11222
rect 16592 10198 16620 15914
rect 16684 13530 16712 16102
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16776 11830 16804 17614
rect 16868 17202 16896 18226
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16868 16658 16896 17138
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16868 15366 16896 16390
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16960 15026 16988 18022
rect 17052 15094 17080 19314
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 12434 16896 13806
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12434 17080 13194
rect 17144 12986 17172 17478
rect 17236 15994 17264 18566
rect 17328 17746 17356 22066
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17420 20806 17448 21830
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17512 18970 17540 23462
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17512 18766 17540 18906
rect 17500 18760 17552 18766
rect 17552 18708 17632 18714
rect 17500 18702 17632 18708
rect 17512 18686 17632 18702
rect 17696 18698 17724 28970
rect 17788 27538 17816 31214
rect 18800 31142 18828 31282
rect 18788 31136 18840 31142
rect 18788 31078 18840 31084
rect 18800 30598 18828 31078
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 18420 30592 18472 30598
rect 18420 30534 18472 30540
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18340 30054 18368 30534
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18340 28422 18368 29990
rect 18432 29510 18460 30534
rect 18800 30054 18828 30534
rect 18788 30048 18840 30054
rect 18788 29990 18840 29996
rect 18972 29776 19024 29782
rect 18972 29718 19024 29724
rect 18880 29572 18932 29578
rect 18880 29514 18932 29520
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18328 28416 18380 28422
rect 18328 28358 18380 28364
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18340 28014 18368 28358
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17972 27470 18000 27950
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18340 26994 18368 27950
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18340 26382 18368 26930
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 26182
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18432 25838 18460 29446
rect 18788 29028 18840 29034
rect 18788 28970 18840 28976
rect 18696 28620 18748 28626
rect 18696 28562 18748 28568
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18524 27878 18552 28018
rect 18616 27878 18644 28086
rect 18512 27872 18564 27878
rect 18510 27840 18512 27849
rect 18604 27872 18656 27878
rect 18564 27840 18566 27849
rect 18604 27814 18656 27820
rect 18510 27775 18566 27784
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 18340 25294 18368 25638
rect 18616 25430 18644 27814
rect 18708 26790 18736 28562
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18604 25424 18656 25430
rect 18604 25366 18656 25372
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18340 25158 18368 25230
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18340 24818 18368 25094
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18432 24614 18460 24686
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17880 22982 17908 23802
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18156 23118 18184 23462
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17880 22166 17908 22918
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17328 16454 17356 17274
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17314 16280 17370 16289
rect 17314 16215 17370 16224
rect 17328 16182 17356 16215
rect 17316 16176 17368 16182
rect 17368 16136 17448 16164
rect 17316 16118 17368 16124
rect 17236 15966 17356 15994
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15337 17264 15846
rect 17328 15706 17356 15966
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17222 15328 17278 15337
rect 17222 15263 17278 15272
rect 17420 15162 17448 16136
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17236 12617 17264 12786
rect 17222 12608 17278 12617
rect 17222 12543 17278 12552
rect 16868 12406 16988 12434
rect 17052 12406 17172 12434
rect 16960 12170 16988 12406
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16684 11082 16712 11766
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16684 9654 16712 11018
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16592 7206 16620 9386
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 9178 16712 9318
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 15948 4542 16068 4570
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 15856 800 15884 2926
rect 15948 2854 15976 4542
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16040 2922 16068 4014
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 16132 2582 16160 6190
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16224 800 16252 4014
rect 16316 2378 16344 6870
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 4554 16436 5510
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16408 4214 16436 4490
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16408 2774 16436 4150
rect 16500 3398 16528 6666
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16408 2746 16528 2774
rect 16500 2650 16528 2746
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16592 800 16620 3062
rect 16776 2446 16804 9862
rect 16868 7546 16896 10610
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16960 7478 16988 9590
rect 17052 9450 17080 11222
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17052 8945 17080 9046
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16868 4826 16896 5850
rect 16960 5234 16988 7142
rect 17052 6730 17080 8366
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17052 4826 17080 5102
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17144 3058 17172 12406
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17236 7886 17264 11698
rect 17328 11286 17356 13670
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17420 13326 17448 13466
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17420 11218 17448 12106
rect 17512 11898 17540 18566
rect 17604 17678 17632 18686
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17592 16992 17644 16998
rect 17696 16980 17724 17682
rect 17788 17542 17816 20878
rect 17880 20398 17908 21830
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17880 19922 17908 20334
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 18340 19854 18368 24550
rect 18432 23526 18460 24550
rect 18524 24206 18552 25094
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23798 18552 24006
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18432 20602 18460 23122
rect 18616 23118 18644 24822
rect 18708 24274 18736 26726
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18512 23044 18564 23050
rect 18512 22986 18564 22992
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 17866 17912 17922 17921
rect 17866 17847 17868 17856
rect 17920 17847 17922 17856
rect 17868 17818 17920 17824
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17880 17270 17908 17818
rect 18340 17746 18368 18022
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17644 16952 17724 16980
rect 17592 16934 17644 16940
rect 17604 13734 17632 16934
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15348 18000 16050
rect 18340 15434 18368 17682
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 17880 15320 18000 15348
rect 17880 15144 17908 15320
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17880 15116 18368 15144
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17604 12986 17632 13466
rect 18340 13326 18368 15116
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17328 9586 17356 11018
rect 17420 9722 17448 11154
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17420 8838 17448 9318
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17314 8528 17370 8537
rect 17314 8463 17316 8472
rect 17368 8463 17370 8472
rect 17316 8434 17368 8440
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17420 7002 17448 7210
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17314 6896 17370 6905
rect 17314 6831 17370 6840
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 4486 17264 6258
rect 17328 5817 17356 6831
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17314 5808 17370 5817
rect 17314 5743 17370 5752
rect 17420 5030 17448 6190
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16960 800 16988 2382
rect 17328 800 17356 4490
rect 17512 3534 17540 10474
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17604 3194 17632 11766
rect 17880 11354 17908 11834
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17682 10704 17738 10713
rect 17682 10639 17684 10648
rect 17736 10639 17738 10648
rect 17776 10668 17828 10674
rect 17684 10610 17736 10616
rect 17776 10610 17828 10616
rect 17682 10568 17738 10577
rect 17682 10503 17738 10512
rect 17696 10062 17724 10503
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17696 7954 17724 8978
rect 17788 8022 17816 10610
rect 17880 9994 17908 11290
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10742 18368 12786
rect 18432 12617 18460 17478
rect 18524 17270 18552 22986
rect 18616 22778 18644 23054
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18616 22506 18644 22714
rect 18708 22642 18736 22918
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18604 22500 18656 22506
rect 18604 22442 18656 22448
rect 18708 22234 18736 22578
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18694 22128 18750 22137
rect 18694 22063 18750 22072
rect 18708 21690 18736 22063
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18708 21434 18736 21626
rect 18800 21622 18828 28970
rect 18892 28762 18920 29514
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18984 25974 19012 29718
rect 19076 29102 19104 32166
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19168 29306 19196 29446
rect 19260 29306 19288 35498
rect 19996 35018 20024 44950
rect 20720 43784 20772 43790
rect 20720 43726 20772 43732
rect 20536 35556 20588 35562
rect 20536 35498 20588 35504
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 20260 35012 20312 35018
rect 20260 34954 20312 34960
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19352 32314 19380 33934
rect 19708 33924 19760 33930
rect 19708 33866 19760 33872
rect 20168 33924 20220 33930
rect 20168 33866 20220 33872
rect 19720 33318 19748 33866
rect 20180 33658 20208 33866
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 19708 33312 19760 33318
rect 19708 33254 19760 33260
rect 20076 32496 20128 32502
rect 20180 32450 20208 33594
rect 20128 32444 20208 32450
rect 20076 32438 20208 32444
rect 20088 32422 20208 32438
rect 19352 32286 19472 32314
rect 19444 32230 19472 32286
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19444 31822 19472 32166
rect 20180 32026 20208 32422
rect 20168 32020 20220 32026
rect 20168 31962 20220 31968
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19444 30802 19472 31758
rect 19720 31482 19748 31826
rect 20180 31754 20208 31962
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 19708 31476 19760 31482
rect 19708 31418 19760 31424
rect 20180 31414 20208 31690
rect 20168 31408 20220 31414
rect 20168 31350 20220 31356
rect 20272 31346 20300 34954
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 20260 30592 20312 30598
rect 20260 30534 20312 30540
rect 20272 30394 20300 30534
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19352 29306 19380 29650
rect 19996 29510 20024 30262
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19996 29238 20024 29446
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 19064 29096 19116 29102
rect 19064 29038 19116 29044
rect 19076 28490 19104 29038
rect 19064 28484 19116 28490
rect 19064 28426 19116 28432
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19800 28416 19852 28422
rect 19800 28358 19852 28364
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19444 26382 19472 26726
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 19076 25702 19104 25978
rect 19064 25696 19116 25702
rect 19064 25638 19116 25644
rect 19444 24750 19472 26318
rect 19156 24744 19208 24750
rect 19156 24686 19208 24692
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18708 21406 18828 21434
rect 18800 21350 18828 21406
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18512 17264 18564 17270
rect 18512 17206 18564 17212
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16658 18644 17070
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18524 13802 18552 15642
rect 18616 15570 18644 16594
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18418 12608 18474 12617
rect 18418 12543 18474 12552
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11898 18460 12038
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18418 10160 18474 10169
rect 18418 10095 18420 10104
rect 18472 10095 18474 10104
rect 18420 10066 18472 10072
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 18236 9920 18288 9926
rect 18288 9880 18368 9908
rect 18236 9862 18288 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17972 9042 18000 9114
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17880 8498 17908 8842
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18340 7546 18368 9880
rect 18432 8906 18460 10066
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17880 6730 17908 7414
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17696 5914 17724 6666
rect 17880 6458 17908 6666
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17788 5914 17816 6258
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17682 5400 17738 5409
rect 17950 5403 18258 5412
rect 17682 5335 17738 5344
rect 17696 5030 17724 5335
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17880 4282 17908 5102
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 18340 4078 18368 5510
rect 18432 5166 18460 8434
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18524 4146 18552 13194
rect 18616 11558 18644 14826
rect 18708 12306 18736 19654
rect 18800 19242 18828 21286
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18800 14074 18828 17206
rect 18892 16182 18920 24278
rect 19168 24274 19196 24686
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 18972 24132 19024 24138
rect 18972 24074 19024 24080
rect 18984 23526 19012 24074
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 19062 23488 19118 23497
rect 18984 19281 19012 23462
rect 19062 23423 19118 23432
rect 19076 23186 19104 23423
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 19076 22273 19104 23122
rect 19062 22264 19118 22273
rect 19062 22199 19118 22208
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19076 20874 19104 22034
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 19168 20466 19196 24210
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19260 20942 19288 23734
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18970 19272 19026 19281
rect 18970 19207 19026 19216
rect 19076 16402 19104 20198
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19168 18834 19196 19110
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 18984 16374 19104 16402
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18800 12782 18828 14010
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18786 12608 18842 12617
rect 18786 12543 18842 12552
rect 18800 12442 18828 12543
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18800 11150 18828 12378
rect 18892 11898 18920 14962
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18984 10577 19012 16374
rect 19064 15360 19116 15366
rect 19168 15348 19196 18022
rect 19260 17610 19288 19450
rect 19444 17678 19472 23190
rect 19536 19854 19564 28358
rect 19812 28218 19840 28358
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19708 25220 19760 25226
rect 19708 25162 19760 25168
rect 19720 24993 19748 25162
rect 19706 24984 19762 24993
rect 19904 24954 19932 25366
rect 19706 24919 19762 24928
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19628 22778 19656 23666
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19720 22658 19748 24550
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19628 22630 19748 22658
rect 19628 21894 19656 22630
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19720 21486 19748 22510
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 16182 19380 16458
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19116 15320 19196 15348
rect 19064 15302 19116 15308
rect 19076 14890 19104 15302
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 19076 14074 19104 14826
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19076 13938 19104 14010
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19076 12374 19104 12922
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 19168 12306 19196 12786
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 18970 10568 19026 10577
rect 18970 10503 19026 10512
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18616 7342 18644 10066
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18708 7546 18736 9590
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18616 5166 18644 7278
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17696 800 17724 3538
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18432 2774 18460 4014
rect 18616 2774 18644 4694
rect 18708 4146 18736 6938
rect 18800 6338 18828 10406
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18984 9722 19012 9998
rect 18972 9716 19024 9722
rect 19260 9704 19288 15846
rect 19352 13326 19380 16118
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19352 12238 19380 13262
rect 19432 12436 19484 12442
rect 19536 12434 19564 16390
rect 19628 15434 19656 20946
rect 19720 20346 19748 21422
rect 19812 20890 19840 23530
rect 19904 22094 19932 24890
rect 19996 23662 20024 29174
rect 20088 26058 20116 29990
rect 20364 29714 20392 34682
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20456 30190 20484 33254
rect 20548 30326 20576 35498
rect 20732 34406 20760 43726
rect 20996 42560 21048 42566
rect 20996 42502 21048 42508
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20812 32836 20864 32842
rect 20812 32778 20864 32784
rect 20824 32366 20852 32778
rect 20812 32360 20864 32366
rect 20812 32302 20864 32308
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 20916 30666 20944 31826
rect 20904 30660 20956 30666
rect 20904 30602 20956 30608
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20456 28558 20484 29582
rect 20916 28626 20944 30602
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20456 28014 20484 28494
rect 20812 28144 20864 28150
rect 20812 28086 20864 28092
rect 20444 28008 20496 28014
rect 20444 27950 20496 27956
rect 20456 26926 20484 27950
rect 20824 27402 20852 28086
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 26314 20208 26726
rect 20350 26480 20406 26489
rect 20732 26450 20760 27270
rect 20824 26790 20852 27338
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26518 20852 26726
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20350 26415 20406 26424
rect 20720 26444 20772 26450
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20180 26194 20208 26250
rect 20180 26166 20300 26194
rect 20088 26030 20208 26058
rect 20076 24744 20128 24750
rect 20076 24686 20128 24692
rect 20088 24070 20116 24686
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19996 23497 20024 23598
rect 19982 23488 20038 23497
rect 19982 23423 20038 23432
rect 20088 23186 20116 24006
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19904 22066 20116 22094
rect 20088 21894 20116 22066
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19996 21622 20024 21830
rect 20088 21690 20116 21830
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19812 20862 20024 20890
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 19720 20318 19840 20346
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19720 19417 19748 20198
rect 19812 19786 19840 20318
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19706 19408 19762 19417
rect 19706 19343 19762 19352
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19628 14770 19656 15370
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 14958 19840 15302
rect 19904 15162 19932 20742
rect 19996 16250 20024 20862
rect 20180 20534 20208 26030
rect 20272 24886 20300 26166
rect 20364 25430 20392 26415
rect 20720 26386 20772 26392
rect 20352 25424 20404 25430
rect 20352 25366 20404 25372
rect 20364 25294 20392 25366
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 20260 24880 20312 24886
rect 20260 24822 20312 24828
rect 20272 24562 20300 24822
rect 20272 24534 20392 24562
rect 20364 24138 20392 24534
rect 20352 24132 20404 24138
rect 20444 24132 20496 24138
rect 20404 24092 20444 24120
rect 20352 24074 20404 24080
rect 20444 24074 20496 24080
rect 20732 23798 20760 26386
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 20916 24138 20944 25774
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20272 23118 20300 23734
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20824 23186 20852 23666
rect 20916 23662 20944 24074
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 22438 20484 22578
rect 20812 22500 20864 22506
rect 20812 22442 20864 22448
rect 20444 22432 20496 22438
rect 20442 22400 20444 22409
rect 20720 22432 20772 22438
rect 20496 22400 20498 22409
rect 20720 22374 20772 22380
rect 20442 22335 20498 22344
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19628 14742 19840 14770
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19628 14006 19656 14282
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19536 12406 19748 12434
rect 19432 12378 19484 12384
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19444 11762 19472 12378
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19352 10130 19380 11154
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 18972 9658 19024 9664
rect 19076 9676 19288 9704
rect 19076 9042 19104 9676
rect 19154 9616 19210 9625
rect 19154 9551 19210 9560
rect 19248 9580 19300 9586
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 19168 8974 19196 9551
rect 19248 9522 19300 9528
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18800 6310 18920 6338
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18892 3942 18920 6310
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18340 2746 18460 2774
rect 18524 2746 18644 2774
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 11900 734 12112 762
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 2746
rect 18524 2394 18552 2746
rect 18432 2366 18552 2394
rect 18432 800 18460 2366
rect 18800 800 18828 3402
rect 18892 2650 18920 3470
rect 18984 2774 19012 6394
rect 19076 3670 19104 8366
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19168 6390 19196 6598
rect 19156 6384 19208 6390
rect 19156 6326 19208 6332
rect 19260 3738 19288 9522
rect 19352 9178 19380 10066
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 5778 19380 7686
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19352 2774 19380 5578
rect 18984 2746 19104 2774
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 19076 2446 19104 2746
rect 19168 2746 19380 2774
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19168 800 19196 2746
rect 19444 2446 19472 11494
rect 19616 10736 19668 10742
rect 19720 10724 19748 12406
rect 19812 11830 19840 14742
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19904 12442 19932 14350
rect 19996 12986 20024 16050
rect 20088 15094 20116 19110
rect 20180 17338 20208 19722
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20272 16658 20300 19858
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 16250 20300 16594
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20272 15570 20300 16186
rect 20364 16182 20392 21830
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 19514 20484 21286
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20548 19378 20576 20334
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20456 14770 20484 17002
rect 20640 16658 20668 22034
rect 20732 19514 20760 22374
rect 20824 20534 20852 22442
rect 20916 21894 20944 23598
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 21008 18714 21036 42502
rect 21744 35698 21772 46038
rect 21836 43858 21864 47942
rect 21824 43852 21876 43858
rect 21824 43794 21876 43800
rect 22008 39296 22060 39302
rect 22008 39238 22060 39244
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 21100 35601 21128 35634
rect 21272 35624 21324 35630
rect 21086 35592 21142 35601
rect 21272 35566 21324 35572
rect 21086 35527 21142 35536
rect 21284 33946 21312 35566
rect 21744 35290 21772 35634
rect 21732 35284 21784 35290
rect 21732 35226 21784 35232
rect 21192 33918 21312 33946
rect 21192 33862 21220 33918
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21192 32502 21220 33798
rect 21180 32496 21232 32502
rect 21180 32438 21232 32444
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 21100 32026 21128 32166
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 21284 28082 21312 29106
rect 21364 28620 21416 28626
rect 21364 28562 21416 28568
rect 21376 28490 21404 28562
rect 21364 28484 21416 28490
rect 21364 28426 21416 28432
rect 21376 28150 21404 28426
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21284 27946 21312 28018
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21272 26852 21324 26858
rect 21272 26794 21324 26800
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 21100 21146 21128 22170
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 21100 20398 21128 21082
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 20824 18686 21036 18714
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20548 15366 20576 16594
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20364 14742 20484 14770
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20180 13938 20208 14214
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19668 10696 19748 10724
rect 19616 10678 19668 10684
rect 19616 10600 19668 10606
rect 19614 10568 19616 10577
rect 19668 10568 19670 10577
rect 19614 10503 19670 10512
rect 19524 9920 19576 9926
rect 19576 9880 19656 9908
rect 19524 9862 19576 9868
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19536 3534 19564 8842
rect 19628 4622 19656 9880
rect 19720 5778 19748 10696
rect 19812 9926 19840 10950
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19812 9450 19840 9590
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19812 8906 19840 9386
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19812 7750 19840 8842
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7546 19840 7686
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19812 6934 19840 7482
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19812 5302 19840 6870
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19812 4214 19840 5238
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19904 3058 19932 12106
rect 20088 11830 20116 13330
rect 20272 12374 20300 14214
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20364 12186 20392 14742
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20180 12158 20392 12186
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 19984 11688 20036 11694
rect 20180 11642 20208 12158
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11898 20392 12038
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 19984 11630 20036 11636
rect 19996 11150 20024 11630
rect 20088 11614 20208 11642
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19996 10810 20024 10950
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19996 10266 20024 10610
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19996 9110 20024 9862
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 20088 7886 20116 11614
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20088 5681 20116 6598
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 20180 3534 20208 11494
rect 20272 11354 20300 11494
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20364 10792 20392 11698
rect 20456 11354 20484 14214
rect 20640 12850 20668 16594
rect 20732 15570 20760 17478
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20732 13190 20760 14554
rect 20824 14550 20852 18686
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20824 13002 20852 14486
rect 20732 12974 20852 13002
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20272 10764 20392 10792
rect 20272 9994 20300 10764
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20456 10441 20484 10542
rect 20442 10432 20498 10441
rect 20442 10367 20498 10376
rect 20548 10282 20576 12310
rect 20640 11778 20668 12650
rect 20732 12306 20760 12974
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20732 11898 20760 12242
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20640 11750 20760 11778
rect 20916 11762 20944 18566
rect 21088 18080 21140 18086
rect 21086 18048 21088 18057
rect 21140 18048 21142 18057
rect 21086 17983 21142 17992
rect 21192 17678 21220 19994
rect 21284 18290 21312 26794
rect 21468 25906 21496 31282
rect 21652 28422 21680 31622
rect 21744 31414 21772 35226
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21836 33930 21864 34342
rect 21824 33924 21876 33930
rect 21824 33866 21876 33872
rect 21836 33658 21864 33866
rect 21824 33652 21876 33658
rect 21824 33594 21876 33600
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21836 32434 21864 32710
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21836 32230 21864 32370
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21548 28144 21600 28150
rect 21548 28086 21600 28092
rect 21560 27878 21588 28086
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21560 27130 21588 27814
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21468 25702 21496 25842
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21376 18170 21404 24550
rect 21468 22642 21496 25638
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21560 25294 21588 25434
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21548 24676 21600 24682
rect 21548 24618 21600 24624
rect 21560 24070 21588 24618
rect 21652 24410 21680 27814
rect 21640 24404 21692 24410
rect 21640 24346 21692 24352
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21560 23798 21588 24006
rect 21548 23792 21600 23798
rect 21548 23734 21600 23740
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21560 22030 21588 23734
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 22710 21680 23054
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21560 21622 21588 21966
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21560 21350 21588 21558
rect 21640 21412 21692 21418
rect 21640 21354 21692 21360
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21560 19786 21588 21286
rect 21652 20534 21680 21354
rect 21744 20602 21772 29990
rect 21836 29170 21864 32166
rect 22020 31890 22048 39238
rect 22112 35894 22140 53926
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53650 23336 55186
rect 23296 53644 23348 53650
rect 23296 53586 23348 53592
rect 22560 53576 22612 53582
rect 22560 53518 22612 53524
rect 22572 53242 22600 53518
rect 22744 53508 22796 53514
rect 22744 53450 22796 53456
rect 22652 53440 22704 53446
rect 22652 53382 22704 53388
rect 22560 53236 22612 53242
rect 22560 53178 22612 53184
rect 22112 35866 22416 35894
rect 22284 35148 22336 35154
rect 22284 35090 22336 35096
rect 22192 34400 22244 34406
rect 22192 34342 22244 34348
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22112 33318 22140 34138
rect 22100 33312 22152 33318
rect 22100 33254 22152 33260
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31414 22048 31622
rect 22008 31408 22060 31414
rect 22008 31350 22060 31356
rect 22112 29850 22140 32166
rect 22204 30326 22232 34342
rect 22296 33590 22324 35090
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22296 33114 22324 33526
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 22388 31754 22416 35866
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 22572 34202 22600 35566
rect 22664 34406 22692 53382
rect 22756 35894 22784 53450
rect 23308 53242 23336 53586
rect 23400 53582 23428 56063
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 23400 53242 23428 53518
rect 23664 53440 23716 53446
rect 23664 53382 23716 53388
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 23388 53236 23440 53242
rect 23388 53178 23440 53184
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23572 52624 23624 52630
rect 23572 52566 23624 52572
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 23388 43784 23440 43790
rect 23388 43726 23440 43732
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23296 40180 23348 40186
rect 23296 40122 23348 40128
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22756 35866 22876 35894
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22560 34196 22612 34202
rect 22560 34138 22612 34144
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 22664 33810 22692 34002
rect 22572 33782 22692 33810
rect 22572 33658 22600 33782
rect 22560 33652 22612 33658
rect 22560 33594 22612 33600
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22296 31726 22416 31754
rect 22192 30320 22244 30326
rect 22192 30262 22244 30268
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21916 28688 21968 28694
rect 21916 28630 21968 28636
rect 21928 23866 21956 28630
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22112 27674 22140 28562
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22100 27668 22152 27674
rect 22100 27610 22152 27616
rect 22008 27396 22060 27402
rect 22008 27338 22060 27344
rect 22020 26790 22048 27338
rect 22100 27056 22152 27062
rect 22100 26998 22152 27004
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 22112 26586 22140 26998
rect 22204 26994 22232 28358
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22296 26602 22324 31726
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22388 31226 22416 31622
rect 22480 31346 22508 32370
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 22388 31198 22508 31226
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 22388 30802 22416 31078
rect 22376 30796 22428 30802
rect 22376 30738 22428 30744
rect 22376 30660 22428 30666
rect 22376 30602 22428 30608
rect 22388 27130 22416 30602
rect 22480 30036 22508 31198
rect 22572 30190 22600 33594
rect 22650 33144 22706 33153
rect 22650 33079 22706 33088
rect 22664 31686 22692 33079
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22664 30938 22692 31350
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22652 30796 22704 30802
rect 22652 30738 22704 30744
rect 22560 30184 22612 30190
rect 22560 30126 22612 30132
rect 22480 30008 22600 30036
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22204 26574 22324 26602
rect 22204 26042 22232 26574
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 22094 21956 23462
rect 22020 23050 22048 25638
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22204 23730 22232 25094
rect 22296 24750 22324 26386
rect 22388 26314 22416 26930
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22480 26042 22508 29446
rect 22572 28150 22600 30008
rect 22664 28422 22692 30738
rect 22756 30326 22784 34886
rect 22848 32230 22876 35866
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23204 33924 23256 33930
rect 23204 33866 23256 33872
rect 23216 33402 23244 33866
rect 23308 33538 23336 40122
rect 23400 34066 23428 43726
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23308 33510 23428 33538
rect 23296 33448 23348 33454
rect 23216 33396 23296 33402
rect 23216 33390 23348 33396
rect 23216 33374 23336 33390
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23308 32978 23336 33374
rect 23296 32972 23348 32978
rect 23296 32914 23348 32920
rect 23204 32836 23256 32842
rect 23204 32778 23256 32784
rect 23216 32502 23244 32778
rect 23204 32496 23256 32502
rect 23204 32438 23256 32444
rect 23308 32434 23336 32914
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22836 31952 22888 31958
rect 22836 31894 22888 31900
rect 22744 30320 22796 30326
rect 22744 30262 22796 30268
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22560 28144 22612 28150
rect 22560 28086 22612 28092
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 27062 22600 27950
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22296 24138 22324 24686
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 22642 22140 22918
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 21928 22066 22048 22094
rect 22020 21894 22048 22066
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22572 21690 22600 26454
rect 22664 24818 22692 27270
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22756 24750 22784 27814
rect 22848 27130 22876 31894
rect 23400 31890 23428 33510
rect 23584 33114 23612 52566
rect 23572 33108 23624 33114
rect 23572 33050 23624 33056
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23032 31414 23060 31758
rect 23676 31754 23704 53382
rect 23848 52896 23900 52902
rect 23848 52838 23900 52844
rect 24124 52896 24176 52902
rect 24124 52838 24176 52844
rect 23860 32570 23888 52838
rect 23848 32564 23900 32570
rect 23848 32506 23900 32512
rect 23756 32496 23808 32502
rect 23808 32444 23888 32450
rect 23756 32438 23888 32444
rect 23768 32422 23888 32438
rect 23584 31726 23704 31754
rect 23860 31754 23888 32422
rect 23860 31726 24072 31754
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23308 29102 23336 30126
rect 23388 29776 23440 29782
rect 23388 29718 23440 29724
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 22940 28150 22968 28630
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 23400 27962 23428 29718
rect 23584 29306 23612 31726
rect 24044 31686 24072 31726
rect 24032 31680 24084 31686
rect 24032 31622 24084 31628
rect 24044 31346 24072 31622
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 23756 31136 23808 31142
rect 23676 31084 23756 31090
rect 23676 31078 23808 31084
rect 23676 31062 23796 31078
rect 23676 30190 23704 31062
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 23492 28914 23520 29038
rect 23492 28886 23612 28914
rect 23308 27934 23428 27962
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23308 26382 23336 27934
rect 23584 27878 23612 28886
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23400 27674 23428 27814
rect 23388 27668 23440 27674
rect 23388 27610 23440 27616
rect 23584 27538 23612 27814
rect 23572 27532 23624 27538
rect 23572 27474 23624 27480
rect 23584 26926 23612 27474
rect 23676 27130 23704 30126
rect 24032 29504 24084 29510
rect 24032 29446 24084 29452
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23768 28762 23796 29038
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 23296 24744 23348 24750
rect 23296 24686 23348 24692
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24342 23336 24686
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 23204 23656 23256 23662
rect 23308 23610 23336 24278
rect 23256 23604 23336 23610
rect 23204 23598 23336 23604
rect 23216 23582 23336 23598
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 22001 22876 22510
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22030 23336 23582
rect 23296 22024 23348 22030
rect 22834 21992 22890 22001
rect 23296 21966 23348 21972
rect 22834 21927 22890 21936
rect 23020 21956 23072 21962
rect 23020 21898 23072 21904
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 19310 21680 19654
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21284 18142 21404 18170
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21008 16522 21036 17206
rect 21284 16794 21312 18142
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15706 21496 15846
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21284 15026 21312 15370
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21744 14482 21772 20198
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21836 17270 21864 19110
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21928 16697 21956 17614
rect 21914 16688 21970 16697
rect 21914 16623 21970 16632
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 12782 21036 13670
rect 21192 13462 21220 14010
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21100 12850 21128 13398
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 21284 12434 21312 13806
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21192 12406 21312 12434
rect 21364 12436 21416 12442
rect 20732 11354 20760 11750
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20640 10606 20668 11222
rect 20732 11150 20760 11290
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20456 10254 20576 10282
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 20352 8832 20404 8838
rect 20456 8820 20484 10254
rect 20536 10192 20588 10198
rect 20588 10140 20760 10146
rect 20536 10134 20760 10140
rect 20548 10118 20760 10134
rect 20732 9654 20760 10118
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20404 8792 20484 8820
rect 20352 8774 20404 8780
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20272 5302 20300 6326
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20260 4004 20312 4010
rect 20260 3946 20312 3952
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19536 800 19564 2382
rect 19904 800 19932 2790
rect 20272 800 20300 3946
rect 20364 3738 20392 8774
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20456 2650 20484 8366
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20640 7546 20668 8298
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20548 5234 20576 7414
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6458 20668 6598
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20824 5710 20852 11018
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 9722 20944 10066
rect 21100 9722 21128 10610
rect 21192 9874 21220 12406
rect 21468 12434 21496 12582
rect 21468 12406 21588 12434
rect 21364 12378 21416 12384
rect 21376 12322 21404 12378
rect 21272 12300 21324 12306
rect 21376 12294 21496 12322
rect 21272 12242 21324 12248
rect 21284 10606 21312 12242
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21376 10130 21404 12106
rect 21468 12073 21496 12294
rect 21454 12064 21510 12073
rect 21454 11999 21510 12008
rect 21468 11898 21496 11999
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21468 11150 21496 11562
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21468 10606 21496 10950
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21560 10130 21588 12406
rect 21836 11558 21864 15098
rect 22020 14550 22048 21286
rect 22204 21010 22232 21490
rect 22836 21412 22888 21418
rect 22836 21354 22888 21360
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22112 15570 22140 19382
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 18290 22232 18566
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 17338 22232 17614
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22296 16794 22324 17206
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22284 16788 22336 16794
rect 22204 16748 22284 16776
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22204 15434 22232 16748
rect 22284 16730 22336 16736
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22296 16182 22324 16526
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22008 14544 22060 14550
rect 22008 14486 22060 14492
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21376 9994 21404 10066
rect 21364 9988 21416 9994
rect 21416 9948 21588 9976
rect 21364 9930 21416 9936
rect 21192 9846 21404 9874
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21376 9382 21404 9846
rect 21560 9654 21588 9948
rect 21652 9926 21680 10474
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21008 7290 21036 8978
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8634 21220 8842
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21100 7410 21128 7754
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21284 7342 21312 8774
rect 21272 7336 21324 7342
rect 21008 7262 21128 7290
rect 21272 7278 21324 7284
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20548 4690 20576 5170
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4214 20576 4490
rect 20536 4208 20588 4214
rect 20536 4150 20588 4156
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20548 2038 20576 3878
rect 20732 2774 20760 5578
rect 20916 5137 20944 7142
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20902 5128 20958 5137
rect 20902 5063 20958 5072
rect 21008 4146 21036 6666
rect 21100 5302 21128 7262
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21088 5296 21140 5302
rect 21088 5238 21140 5244
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21100 4486 21128 5102
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20640 2746 20760 2774
rect 20536 2032 20588 2038
rect 20536 1974 20588 1980
rect 20640 800 20668 2746
rect 20916 2514 20944 4082
rect 21100 4078 21128 4422
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 21008 800 21036 3334
rect 21100 3194 21128 3334
rect 21192 3194 21220 7210
rect 21284 6798 21312 7278
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21270 5672 21326 5681
rect 21270 5607 21326 5616
rect 21284 5302 21312 5607
rect 21272 5296 21324 5302
rect 21272 5238 21324 5244
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21284 4010 21312 5102
rect 21376 4486 21404 9318
rect 21468 8974 21496 9590
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21468 6934 21496 8434
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 21560 6730 21588 8298
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21652 6458 21680 6802
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21468 5914 21496 6258
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21468 4214 21496 5170
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21376 800 21404 2926
rect 21560 2774 21588 6326
rect 21652 4554 21680 6394
rect 21744 6118 21772 10950
rect 21836 8362 21864 11494
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21928 8106 21956 13262
rect 22020 12986 22048 13874
rect 22112 12986 22140 14962
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22204 13190 22232 13806
rect 22296 13734 22324 15506
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22204 12850 22232 13126
rect 22388 12918 22416 16934
rect 22480 14006 22508 19450
rect 22756 18766 22784 20198
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22572 13138 22600 17478
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 14074 22692 16526
rect 22756 16182 22784 16730
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22756 16046 22784 16118
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22744 15632 22796 15638
rect 22744 15574 22796 15580
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22480 13110 22600 13138
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22112 10538 22140 12786
rect 22204 12238 22232 12786
rect 22480 12594 22508 13110
rect 22296 12566 22508 12594
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22100 10532 22152 10538
rect 22100 10474 22152 10480
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22020 8294 22048 10406
rect 22204 9994 22232 10746
rect 22296 10674 22324 12566
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22468 10464 22520 10470
rect 22466 10432 22468 10441
rect 22520 10432 22522 10441
rect 22466 10367 22522 10376
rect 22572 10062 22600 12310
rect 22664 11218 22692 13670
rect 22756 11286 22784 15574
rect 22848 15094 22876 21354
rect 23032 21350 23060 21898
rect 23308 21690 23336 21966
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 19310 23336 21286
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23216 16998 23244 17750
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23400 16266 23428 25638
rect 23584 24750 23612 26862
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23662 23520 24006
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23492 21486 23520 23598
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23584 20602 23612 21422
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23492 18290 23520 20266
rect 23584 19446 23612 20334
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23676 19446 23704 19994
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23584 17660 23612 19382
rect 23492 17632 23612 17660
rect 23664 17672 23716 17678
rect 23492 17202 23520 17632
rect 23664 17614 23716 17620
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23308 16238 23428 16266
rect 23492 16266 23520 17138
rect 23676 16794 23704 17614
rect 23768 17270 23796 28698
rect 23940 28552 23992 28558
rect 23940 28494 23992 28500
rect 23952 28422 23980 28494
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 23846 27704 23902 27713
rect 23846 27639 23902 27648
rect 23860 26382 23888 27639
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 23860 25430 23888 26318
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23952 25498 23980 25842
rect 23940 25492 23992 25498
rect 23940 25434 23992 25440
rect 23848 25424 23900 25430
rect 23848 25366 23900 25372
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23860 24449 23888 25162
rect 23846 24440 23902 24449
rect 23846 24375 23902 24384
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23860 22234 23888 23054
rect 23952 22642 23980 23462
rect 24044 23118 24072 29446
rect 24136 28014 24164 52838
rect 24504 52698 24532 56200
rect 25318 55448 25374 55457
rect 25318 55383 25374 55392
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24676 53984 24728 53990
rect 24676 53926 24728 53932
rect 24688 53582 24716 53926
rect 24676 53576 24728 53582
rect 24676 53518 24728 53524
rect 24584 53440 24636 53446
rect 24584 53382 24636 53388
rect 24492 52692 24544 52698
rect 24492 52634 24544 52640
rect 24504 52494 24532 52634
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24596 52018 24624 53382
rect 24780 53242 24808 54567
rect 24858 53816 24914 53825
rect 24858 53751 24914 53760
rect 24872 53718 24900 53751
rect 24860 53712 24912 53718
rect 24860 53654 24912 53660
rect 25332 53242 25360 55383
rect 25884 54194 25912 56200
rect 25872 54188 25924 54194
rect 25872 54130 25924 54136
rect 24768 53236 24820 53242
rect 24768 53178 24820 53184
rect 25320 53236 25372 53242
rect 25320 53178 25372 53184
rect 25502 53000 25558 53009
rect 25502 52935 25504 52944
rect 25556 52935 25558 52944
rect 25504 52906 25556 52912
rect 25228 52420 25280 52426
rect 25228 52362 25280 52368
rect 25240 52193 25268 52362
rect 25226 52184 25282 52193
rect 25226 52119 25228 52128
rect 25280 52119 25282 52128
rect 25228 52090 25280 52096
rect 25516 52018 25544 52906
rect 24584 52012 24636 52018
rect 24584 51954 24636 51960
rect 25504 52012 25556 52018
rect 25504 51954 25556 51960
rect 24400 51808 24452 51814
rect 24400 51750 24452 51756
rect 26884 51808 26936 51814
rect 26884 51750 26936 51756
rect 24412 48142 24440 51750
rect 25226 51368 25282 51377
rect 25226 51303 25228 51312
rect 25280 51303 25282 51312
rect 25228 51274 25280 51280
rect 26516 51264 26568 51270
rect 26516 51206 26568 51212
rect 25228 50924 25280 50930
rect 25228 50866 25280 50872
rect 25240 50561 25268 50866
rect 26240 50720 26292 50726
rect 26240 50662 26292 50668
rect 25226 50552 25282 50561
rect 25226 50487 25282 50496
rect 25320 50176 25372 50182
rect 25320 50118 25372 50124
rect 25332 49774 25360 50118
rect 25136 49768 25188 49774
rect 25320 49768 25372 49774
rect 25136 49710 25188 49716
rect 25318 49736 25320 49745
rect 25372 49736 25374 49745
rect 24400 48136 24452 48142
rect 24400 48078 24452 48084
rect 25044 46368 25096 46374
rect 25044 46310 25096 46316
rect 24952 45824 25004 45830
rect 24952 45766 25004 45772
rect 24308 43172 24360 43178
rect 24308 43114 24360 43120
rect 24216 33856 24268 33862
rect 24216 33798 24268 33804
rect 24228 33318 24256 33798
rect 24216 33312 24268 33318
rect 24216 33254 24268 33260
rect 24228 32502 24256 33254
rect 24216 32496 24268 32502
rect 24216 32438 24268 32444
rect 24216 29028 24268 29034
rect 24216 28970 24268 28976
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 24136 24274 24164 24822
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23860 19786 23888 20538
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23846 19544 23902 19553
rect 24044 19514 24072 22918
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 23846 19479 23902 19488
rect 24032 19508 24084 19514
rect 23860 18834 23888 19479
rect 24032 19450 24084 19456
rect 24136 19446 24164 19722
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 24124 17332 24176 17338
rect 24228 17320 24256 28970
rect 24176 17292 24256 17320
rect 24124 17274 24176 17280
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 23846 17096 23902 17105
rect 23846 17031 23902 17040
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23860 16590 23888 17031
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23492 16250 23612 16266
rect 23492 16244 23624 16250
rect 23492 16238 23572 16244
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15586 23336 16238
rect 23492 15586 23520 16238
rect 23572 16186 23624 16192
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23308 15558 23428 15586
rect 23492 15570 23704 15586
rect 23492 15564 23716 15570
rect 23492 15558 23664 15564
rect 23294 15464 23350 15473
rect 23294 15399 23350 15408
rect 23308 15094 23336 15399
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22848 12374 22876 14826
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23204 13864 23256 13870
rect 23308 13818 23336 14350
rect 23400 14346 23428 15558
rect 23664 15506 23716 15512
rect 23768 15434 23796 15846
rect 23756 15428 23808 15434
rect 23756 15370 23808 15376
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 23256 13812 23336 13818
rect 23204 13806 23336 13812
rect 23216 13790 23336 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 12918 23336 13790
rect 23386 13832 23442 13841
rect 23386 13767 23442 13776
rect 23400 13394 23428 13767
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22744 11280 22796 11286
rect 22744 11222 22796 11228
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22848 10606 22876 12174
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11354 23336 11494
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 22836 10600 22888 10606
rect 22650 10568 22706 10577
rect 23308 10577 23336 11154
rect 23400 10742 23428 12582
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 22836 10542 22888 10548
rect 23294 10568 23350 10577
rect 22650 10503 22706 10512
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 22112 9042 22140 9386
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 21928 8078 22048 8106
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21730 5536 21786 5545
rect 21730 5471 21786 5480
rect 21744 4622 21772 5471
rect 21836 4622 21864 7822
rect 22020 6798 22048 8078
rect 22112 7886 22140 8978
rect 22192 8832 22244 8838
rect 22244 8780 22324 8786
rect 22192 8774 22324 8780
rect 22204 8758 22324 8774
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22112 7478 22140 7822
rect 22100 7472 22152 7478
rect 22100 7414 22152 7420
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22204 5522 22232 8434
rect 22296 5710 22324 8758
rect 22388 6905 22416 9862
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22374 6896 22430 6905
rect 22374 6831 22430 6840
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22204 5494 22324 5522
rect 22296 5250 22324 5494
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22204 5222 22324 5250
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22020 3074 22048 4218
rect 22112 3194 22140 5170
rect 22204 3194 22232 5222
rect 22388 4706 22416 6666
rect 22296 4678 22416 4706
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22020 3046 22232 3074
rect 22296 3058 22324 4678
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 21560 2746 21772 2774
rect 21744 800 21772 2746
rect 22204 2666 22232 3046
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22388 2854 22416 4490
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22204 2638 22324 2666
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 22098 2408 22154 2417
rect 22098 2343 22154 2352
rect 22112 1902 22140 2343
rect 22100 1896 22152 1902
rect 22100 1838 22152 1844
rect 22204 1601 22232 2518
rect 22190 1592 22246 1601
rect 22190 1527 22246 1536
rect 22296 1442 22324 2638
rect 22112 1414 22324 1442
rect 22112 800 22140 1414
rect 22480 800 22508 8366
rect 22572 7834 22600 9522
rect 22664 9518 22692 10503
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 9654 22784 10406
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22664 8514 22692 9454
rect 22848 9450 22876 10542
rect 23294 10503 23350 10512
rect 23492 10470 23520 12922
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23400 9722 23520 9738
rect 23388 9716 23520 9722
rect 23440 9710 23520 9716
rect 23388 9658 23440 9664
rect 23492 9654 23520 9710
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23388 8832 23440 8838
rect 23492 8820 23520 9590
rect 23440 8792 23520 8820
rect 23388 8774 23440 8780
rect 22664 8486 22876 8514
rect 22848 7954 22876 8486
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22836 7948 22888 7954
rect 22836 7890 22888 7896
rect 23400 7886 23428 8774
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23388 7880 23440 7886
rect 22572 7806 22692 7834
rect 23388 7822 23440 7828
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22572 2774 22600 7686
rect 22664 7562 22692 7806
rect 22664 7534 22784 7562
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 5030 22692 6734
rect 22756 5574 22784 7534
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6928 22888 6934
rect 22836 6870 22888 6876
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22756 3126 22784 5306
rect 22848 3194 22876 6870
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23308 5681 23336 6802
rect 23400 6390 23428 7414
rect 23492 6934 23520 7958
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23480 6928 23532 6934
rect 23480 6870 23532 6876
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23492 6254 23520 6870
rect 23676 6769 23704 7754
rect 23860 7410 23888 16050
rect 23952 14550 23980 16934
rect 24044 16046 24072 17206
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24044 15620 24072 15982
rect 24124 15632 24176 15638
rect 24044 15592 24124 15620
rect 24176 15592 24256 15620
rect 24124 15574 24176 15580
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 23940 14544 23992 14550
rect 23940 14486 23992 14492
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23662 6760 23718 6769
rect 23662 6695 23718 6704
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23294 5672 23350 5681
rect 23294 5607 23350 5616
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23308 3890 23336 5510
rect 23400 4865 23428 6190
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23768 5794 23796 5850
rect 23768 5766 23888 5794
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23768 5234 23796 5578
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23572 5160 23624 5166
rect 23572 5102 23624 5108
rect 23386 4856 23442 4865
rect 23386 4791 23442 4800
rect 23386 3904 23442 3913
rect 23308 3862 23386 3890
rect 22950 3836 23258 3845
rect 23386 3839 23442 3848
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 22940 3126 22968 3674
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23296 3528 23348 3534
rect 23294 3496 23296 3505
rect 23348 3496 23350 3505
rect 23294 3431 23350 3440
rect 23400 3233 23428 3606
rect 23386 3224 23442 3233
rect 23386 3159 23442 3168
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23400 2854 23428 2994
rect 23584 2990 23612 5102
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23768 4554 23796 4762
rect 23756 4548 23808 4554
rect 23756 4490 23808 4496
rect 23664 4480 23716 4486
rect 23860 4434 23888 5766
rect 23952 5710 23980 14214
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 24044 13326 24072 14010
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24136 12442 24164 14962
rect 24228 13938 24256 15592
rect 24320 14618 24348 43114
rect 24860 41540 24912 41546
rect 24860 41482 24912 41488
rect 24872 41449 24900 41482
rect 24858 41440 24914 41449
rect 24858 41375 24914 41384
rect 24860 40928 24912 40934
rect 24860 40870 24912 40876
rect 24872 35766 24900 40870
rect 24964 40746 24992 45766
rect 25056 40934 25084 46310
rect 25044 40928 25096 40934
rect 25044 40870 25096 40876
rect 24964 40718 25084 40746
rect 24952 40384 25004 40390
rect 24952 40326 25004 40332
rect 24860 35760 24912 35766
rect 24860 35702 24912 35708
rect 24964 35086 24992 40326
rect 25056 35834 25084 40718
rect 25044 35828 25096 35834
rect 25044 35770 25096 35776
rect 24952 35080 25004 35086
rect 24952 35022 25004 35028
rect 24584 33312 24636 33318
rect 24584 33254 24636 33260
rect 24768 33312 24820 33318
rect 24768 33254 24820 33260
rect 24596 32774 24624 33254
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24596 29850 24624 32710
rect 24780 32609 24808 33254
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24766 32600 24822 32609
rect 24766 32535 24822 32544
rect 24964 32366 24992 32914
rect 24952 32360 25004 32366
rect 24872 32308 24952 32314
rect 24872 32302 25004 32308
rect 24872 32286 24992 32302
rect 24676 31136 24728 31142
rect 24676 31078 24728 31084
rect 24688 30598 24716 31078
rect 24676 30592 24728 30598
rect 24676 30534 24728 30540
rect 24688 30258 24716 30534
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29510 24532 29582
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 24504 28529 24532 29446
rect 24596 29306 24624 29786
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24490 28520 24546 28529
rect 24490 28455 24546 28464
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24412 28150 24440 28358
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21486 24440 21830
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24504 18698 24532 28358
rect 24688 28150 24716 30194
rect 24872 30190 24900 32286
rect 25148 32178 25176 49710
rect 25318 49671 25374 49680
rect 25228 49156 25280 49162
rect 25228 49098 25280 49104
rect 25240 48929 25268 49098
rect 25596 49088 25648 49094
rect 25596 49030 25648 49036
rect 25226 48920 25282 48929
rect 25226 48855 25282 48864
rect 25228 48544 25280 48550
rect 25228 48486 25280 48492
rect 25240 48142 25268 48486
rect 25228 48136 25280 48142
rect 25226 48104 25228 48113
rect 25280 48104 25282 48113
rect 25226 48039 25282 48048
rect 25320 47660 25372 47666
rect 25320 47602 25372 47608
rect 25332 47297 25360 47602
rect 25412 47456 25464 47462
rect 25412 47398 25464 47404
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25332 46578 25360 46854
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25320 45280 25372 45286
rect 25320 45222 25372 45228
rect 25332 44878 25360 45222
rect 25320 44872 25372 44878
rect 25318 44840 25320 44849
rect 25372 44840 25374 44849
rect 25318 44775 25374 44784
rect 25320 44736 25372 44742
rect 25320 44678 25372 44684
rect 25228 44396 25280 44402
rect 25228 44338 25280 44344
rect 25240 44033 25268 44338
rect 25226 44024 25282 44033
rect 25226 43959 25282 43968
rect 25228 43648 25280 43654
rect 25228 43590 25280 43596
rect 25240 43314 25268 43590
rect 25228 43308 25280 43314
rect 25228 43250 25280 43256
rect 25240 43217 25268 43250
rect 25226 43208 25282 43217
rect 25226 43143 25282 43152
rect 25228 42628 25280 42634
rect 25228 42570 25280 42576
rect 25240 42401 25268 42570
rect 25226 42392 25282 42401
rect 25226 42327 25282 42336
rect 25228 42016 25280 42022
rect 25228 41958 25280 41964
rect 25240 41614 25268 41958
rect 25228 41608 25280 41614
rect 25226 41576 25228 41585
rect 25280 41576 25282 41585
rect 25226 41511 25282 41520
rect 25332 41290 25360 44678
rect 25240 41262 25360 41290
rect 25240 40390 25268 41262
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25228 40384 25280 40390
rect 25228 40326 25280 40332
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 39137 25360 39374
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25332 38350 25360 38694
rect 25320 38344 25372 38350
rect 25318 38312 25320 38321
rect 25372 38312 25374 38321
rect 25318 38247 25374 38256
rect 25228 37868 25280 37874
rect 25228 37810 25280 37816
rect 25240 37505 25268 37810
rect 25226 37496 25282 37505
rect 25226 37431 25282 37440
rect 25228 37120 25280 37126
rect 25228 37062 25280 37068
rect 25240 36786 25268 37062
rect 25228 36780 25280 36786
rect 25228 36722 25280 36728
rect 25240 36689 25268 36722
rect 25226 36680 25282 36689
rect 25226 36615 25282 36624
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25332 35873 25360 36110
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25332 35086 25360 35430
rect 25320 35080 25372 35086
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25318 34983 25374 34992
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25374 34176
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25332 33425 25360 33934
rect 25318 33416 25374 33425
rect 25424 33386 25452 47398
rect 25504 40384 25556 40390
rect 25504 40326 25556 40332
rect 25516 40118 25544 40326
rect 25504 40112 25556 40118
rect 25504 40054 25556 40060
rect 25516 39953 25544 40054
rect 25502 39944 25558 39953
rect 25502 39879 25558 39888
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25318 33351 25374 33360
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 25412 32836 25464 32842
rect 25412 32778 25464 32784
rect 25228 32768 25280 32774
rect 25228 32710 25280 32716
rect 24964 32150 25176 32178
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24872 29345 24900 29514
rect 24858 29336 24914 29345
rect 24858 29271 24914 29280
rect 24964 29238 24992 32150
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24964 28558 24992 29038
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24952 28144 25004 28150
rect 24952 28086 25004 28092
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24688 27606 24716 27950
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24688 27130 24716 27542
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 24872 26194 24900 27406
rect 24964 26994 24992 28086
rect 25056 27538 25084 31894
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24780 26166 24900 26194
rect 24780 26042 24808 26166
rect 24858 26072 24914 26081
rect 24768 26036 24820 26042
rect 24858 26007 24914 26016
rect 24768 25978 24820 25984
rect 24872 25974 24900 26007
rect 24860 25968 24912 25974
rect 24860 25910 24912 25916
rect 24872 25498 24900 25910
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24676 25424 24728 25430
rect 24676 25366 24728 25372
rect 24688 22778 24716 25366
rect 24964 24970 24992 26522
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 24872 24942 24992 24970
rect 24872 23746 24900 24942
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24964 24410 24992 24754
rect 25056 24750 25084 26386
rect 25148 26314 25176 31078
rect 25240 28558 25268 32710
rect 25424 32230 25452 32778
rect 25412 32224 25464 32230
rect 25412 32166 25464 32172
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25424 28626 25452 32166
rect 25516 31482 25544 38150
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25516 30977 25544 31282
rect 25502 30968 25558 30977
rect 25502 30903 25504 30912
rect 25556 30903 25558 30912
rect 25504 30874 25556 30880
rect 25504 29232 25556 29238
rect 25504 29174 25556 29180
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 25228 28552 25280 28558
rect 25228 28494 25280 28500
rect 25412 27872 25464 27878
rect 25412 27814 25464 27820
rect 25424 27470 25452 27814
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25412 26920 25464 26926
rect 25318 26888 25374 26897
rect 25412 26862 25464 26868
rect 25318 26823 25374 26832
rect 25228 26512 25280 26518
rect 25228 26454 25280 26460
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25056 23866 25084 24686
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 25148 23798 25176 24346
rect 25136 23792 25188 23798
rect 24872 23718 25084 23746
rect 25136 23734 25188 23740
rect 24766 23624 24822 23633
rect 24766 23559 24822 23568
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24780 22574 24808 23559
rect 24860 23180 24912 23186
rect 24860 23122 24912 23128
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24872 22817 24900 23122
rect 24858 22808 24914 22817
rect 24858 22743 24914 22752
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24964 21350 24992 23122
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24582 20360 24638 20369
rect 24582 20295 24638 20304
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24596 18222 24624 20295
rect 24688 20058 24716 20946
rect 24872 20942 24900 21111
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24964 20806 24992 20946
rect 25056 20942 25084 23718
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25148 23050 25176 23462
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 25240 22030 25268 26454
rect 25332 25294 25360 26823
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25332 24410 25360 25230
rect 25424 24750 25452 26862
rect 25516 26489 25544 29174
rect 25502 26480 25558 26489
rect 25502 26415 25558 26424
rect 25608 25770 25636 49030
rect 25872 48000 25924 48006
rect 25872 47942 25924 47948
rect 25688 44192 25740 44198
rect 25688 44134 25740 44140
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 25424 22234 25452 24686
rect 25516 23526 25544 25094
rect 25608 24834 25636 25434
rect 25700 24970 25728 44134
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25792 25498 25820 36518
rect 25884 29034 25912 47942
rect 25964 37664 26016 37670
rect 25964 37606 26016 37612
rect 25872 29028 25924 29034
rect 25872 28970 25924 28976
rect 25872 28688 25924 28694
rect 25872 28630 25924 28636
rect 25884 26246 25912 28630
rect 25872 26240 25924 26246
rect 25872 26182 25924 26188
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25884 25158 25912 26182
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25700 24942 25912 24970
rect 25608 24806 25820 24834
rect 25504 23520 25556 23526
rect 25504 23462 25556 23468
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25516 22094 25544 23258
rect 25424 22066 25544 22094
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24964 19718 24992 20742
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24858 18728 24914 18737
rect 24858 18663 24914 18672
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24688 18057 24716 18566
rect 24872 18358 24900 18663
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24674 18048 24730 18057
rect 24674 17983 24730 17992
rect 24858 17912 24914 17921
rect 24858 17847 24860 17856
rect 24912 17847 24914 17856
rect 24860 17818 24912 17824
rect 24964 17626 24992 19654
rect 25056 17746 25084 20742
rect 25332 20602 25360 21422
rect 25424 21010 25452 22066
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 19514 25176 20334
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25148 17746 25176 19450
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24400 17604 24452 17610
rect 24964 17598 25084 17626
rect 24400 17546 24452 17552
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24412 13938 24440 17546
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24216 13932 24268 13938
rect 24400 13932 24452 13938
rect 24268 13892 24348 13920
rect 24216 13874 24268 13880
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24044 11354 24072 12174
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24044 8022 24072 11086
rect 24136 10810 24164 12174
rect 24124 10804 24176 10810
rect 24124 10746 24176 10752
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 24136 10130 24164 10406
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24136 9654 24164 10066
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24228 8974 24256 13466
rect 24320 13444 24348 13892
rect 24400 13874 24452 13880
rect 24504 13530 24532 14350
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24320 13416 24440 13444
rect 24412 13258 24440 13416
rect 24308 13252 24360 13258
rect 24308 13194 24360 13200
rect 24400 13252 24452 13258
rect 24400 13194 24452 13200
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24044 6254 24072 7346
rect 24032 6248 24084 6254
rect 24030 6216 24032 6225
rect 24084 6216 24086 6225
rect 24030 6151 24086 6160
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 23664 4422 23716 4428
rect 23572 2984 23624 2990
rect 23676 2961 23704 4422
rect 23768 4406 23888 4434
rect 23572 2926 23624 2932
rect 23662 2952 23718 2961
rect 23480 2916 23532 2922
rect 23662 2887 23718 2896
rect 23480 2858 23532 2864
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 22572 2746 22784 2774
rect 22756 2360 22784 2746
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 22756 2332 22876 2360
rect 22848 800 22876 2332
rect 23216 800 23244 2586
rect 23492 1578 23520 2858
rect 23768 2774 23796 4406
rect 23938 4040 23994 4049
rect 23938 3975 23994 3984
rect 23676 2746 23796 2774
rect 23676 2650 23704 2746
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23492 1550 23612 1578
rect 23584 800 23612 1550
rect 23952 800 23980 3975
rect 24136 3058 24164 8298
rect 24216 6112 24268 6118
rect 24216 6054 24268 6060
rect 24228 5778 24256 6054
rect 24320 5914 24348 13194
rect 24412 12986 24440 13194
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24412 6458 24440 11698
rect 24596 10266 24624 15982
rect 24688 14958 24716 16215
rect 24780 15570 24808 17478
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24858 14648 24914 14657
rect 24858 14583 24914 14592
rect 24872 14482 24900 14583
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24766 13016 24822 13025
rect 24766 12951 24822 12960
rect 24780 11694 24808 12951
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 12209 24900 12242
rect 24858 12200 24914 12209
rect 24858 12135 24914 12144
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24872 11393 24900 11562
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24492 8288 24544 8294
rect 24492 8230 24544 8236
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24308 5908 24360 5914
rect 24308 5850 24360 5856
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24308 4480 24360 4486
rect 24308 4422 24360 4428
rect 24320 4146 24348 4422
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 24228 3738 24256 4082
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 24136 2446 24164 2994
rect 24124 2440 24176 2446
rect 24124 2382 24176 2388
rect 24320 800 24348 4082
rect 24504 2922 24532 8230
rect 24596 3126 24624 9862
rect 24964 9586 24992 15642
rect 25056 10826 25084 17598
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 11762 25176 14214
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25792 11558 25820 24806
rect 25884 18426 25912 24942
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25976 11830 26004 37606
rect 26252 35894 26280 50662
rect 26252 35866 26372 35894
rect 26148 34944 26200 34950
rect 26148 34886 26200 34892
rect 26056 33312 26108 33318
rect 26056 33254 26108 33260
rect 26068 28490 26096 33254
rect 26056 28484 26108 28490
rect 26056 28426 26108 28432
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 26068 26382 26096 27338
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 26068 23322 26096 26318
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 26160 17814 26188 34886
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 26252 28218 26280 33798
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26344 28121 26372 35866
rect 26424 33380 26476 33386
rect 26424 33322 26476 33328
rect 26436 29170 26464 33322
rect 26528 30054 26556 51206
rect 26608 40928 26660 40934
rect 26608 40870 26660 40876
rect 26620 32910 26648 40870
rect 26792 36032 26844 36038
rect 26792 35974 26844 35980
rect 26608 32904 26660 32910
rect 26608 32846 26660 32852
rect 26516 30048 26568 30054
rect 26516 29990 26568 29996
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26330 28112 26386 28121
rect 26330 28047 26386 28056
rect 26436 23254 26464 28970
rect 26424 23248 26476 23254
rect 26424 23190 26476 23196
rect 26804 18970 26832 35974
rect 26896 28966 26924 51750
rect 26884 28960 26936 28966
rect 26884 28902 26936 28908
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26148 17808 26200 17814
rect 26148 17750 26200 17756
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25056 10798 25452 10826
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24688 6458 24716 7686
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24780 5710 24808 8774
rect 24872 7426 24900 9318
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 24872 7398 24992 7426
rect 24860 7336 24912 7342
rect 24858 7304 24860 7313
rect 24912 7304 24914 7313
rect 24858 7239 24914 7248
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 24872 6497 24900 6666
rect 24858 6488 24914 6497
rect 24858 6423 24914 6432
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24964 5273 24992 7398
rect 25056 6866 25084 9930
rect 25134 9752 25190 9761
rect 25332 9722 25360 10678
rect 25134 9687 25190 9696
rect 25320 9716 25372 9722
rect 25148 8566 25176 9687
rect 25320 9658 25372 9664
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25320 8084 25372 8090
rect 25148 7478 25176 8055
rect 25320 8026 25372 8032
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25240 6118 25268 6666
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 24950 5264 25006 5273
rect 24950 5199 25006 5208
rect 25240 4593 25268 6054
rect 25226 4584 25282 4593
rect 25226 4519 25282 4528
rect 24766 4040 24822 4049
rect 24766 3975 24822 3984
rect 24780 3126 24808 3975
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 25240 3534 25268 3878
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25056 3194 25084 3470
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 24492 2916 24544 2922
rect 24492 2858 24544 2864
rect 24780 2514 24808 3062
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 25240 2446 25268 3334
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24596 1970 24624 2246
rect 24584 1964 24636 1970
rect 24584 1906 24636 1912
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25332 785 25360 8026
rect 25424 4185 25452 10798
rect 25410 4176 25466 4185
rect 25410 4111 25466 4120
rect 25318 776 25374 785
rect 25318 711 25374 720
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3882 8744 3938 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 5354 9152 5410 9208
rect 4066 6432 4122 6488
rect 5170 3984 5226 4040
rect 5722 3032 5778 3088
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 23386 56072 23442 56128
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7930 3440 7986 3496
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 10230 6160 10286 6216
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 15566 27276 15568 27296
rect 15568 27276 15620 27296
rect 15620 27276 15622 27296
rect 15566 27240 15622 27276
rect 15198 24656 15254 24712
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12070 11600 12126 11656
rect 11150 5072 11206 5128
rect 11150 4528 11206 4584
rect 11242 3984 11298 4040
rect 11794 7964 11796 7984
rect 11796 7964 11848 7984
rect 11848 7964 11850 7984
rect 11794 7928 11850 7964
rect 12438 12416 12494 12472
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12714 12416 12770 12472
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13082 11620 13138 11656
rect 13082 11600 13084 11620
rect 13084 11600 13136 11620
rect 13136 11600 13138 11620
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12254 5752 12310 5808
rect 12254 5344 12310 5400
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13818 13912 13874 13968
rect 12806 8472 12862 8528
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12898 5228 12954 5264
rect 12898 5208 12900 5228
rect 12900 5208 12952 5228
rect 12952 5208 12954 5228
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12806 4020 12808 4040
rect 12808 4020 12860 4040
rect 12860 4020 12862 4040
rect 12806 3984 12862 4020
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13542 8900 13598 8936
rect 13542 8880 13544 8900
rect 13544 8880 13596 8900
rect 13596 8880 13598 8900
rect 14278 12416 14334 12472
rect 14094 10376 14150 10432
rect 13634 6704 13690 6760
rect 13358 3032 13414 3088
rect 14094 6432 14150 6488
rect 13450 2896 13506 2952
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 16118 28056 16174 28112
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 14738 12416 14794 12472
rect 14646 11500 14648 11520
rect 14648 11500 14700 11520
rect 14700 11500 14702 11520
rect 14646 11464 14702 11500
rect 15382 12552 15438 12608
rect 14370 6840 14426 6896
rect 14370 3984 14426 4040
rect 15750 12552 15806 12608
rect 15290 5616 15346 5672
rect 15658 3576 15714 3632
rect 17406 25780 17408 25800
rect 17408 25780 17460 25800
rect 17460 25780 17462 25800
rect 17406 25744 17462 25780
rect 17314 22752 17370 22808
rect 16210 8336 16266 8392
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 18510 27820 18512 27840
rect 18512 27820 18564 27840
rect 18564 27820 18566 27840
rect 18510 27784 18566 27820
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17314 16224 17370 16280
rect 17222 15272 17278 15328
rect 17222 12552 17278 12608
rect 17038 8880 17094 8936
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17866 17876 17922 17912
rect 17866 17856 17868 17876
rect 17868 17856 17920 17876
rect 17920 17856 17922 17876
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17314 8492 17370 8528
rect 17314 8472 17316 8492
rect 17316 8472 17368 8492
rect 17368 8472 17370 8492
rect 17314 6840 17370 6896
rect 17314 5752 17370 5808
rect 17682 10668 17738 10704
rect 17682 10648 17684 10668
rect 17684 10648 17736 10668
rect 17736 10648 17738 10668
rect 17682 10512 17738 10568
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18694 22072 18750 22128
rect 18418 12552 18474 12608
rect 18418 10124 18474 10160
rect 18418 10104 18420 10124
rect 18420 10104 18472 10124
rect 18472 10104 18474 10124
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17682 5344 17738 5400
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19062 23432 19118 23488
rect 19062 22208 19118 22264
rect 18970 19216 19026 19272
rect 18786 12552 18842 12608
rect 19706 24928 19762 24984
rect 18970 10512 19026 10568
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 20350 26424 20406 26480
rect 19982 23432 20038 23488
rect 19706 19352 19762 19408
rect 20442 22380 20444 22400
rect 20444 22380 20496 22400
rect 20496 22380 20498 22400
rect 20442 22344 20498 22380
rect 19154 9560 19210 9616
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21086 35536 21142 35592
rect 19614 10548 19616 10568
rect 19616 10548 19668 10568
rect 19668 10548 19670 10568
rect 19614 10512 19670 10548
rect 20074 5616 20130 5672
rect 20442 10376 20498 10432
rect 21086 18028 21088 18048
rect 21088 18028 21140 18048
rect 21140 18028 21142 18048
rect 21086 17992 21142 18028
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22650 33088 22706 33144
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22834 21936 22890 21992
rect 21914 16632 21970 16688
rect 21454 12008 21510 12064
rect 20902 5072 20958 5128
rect 21270 5616 21326 5672
rect 22466 10412 22468 10432
rect 22468 10412 22520 10432
rect 22520 10412 22522 10432
rect 22466 10376 22522 10412
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23846 27648 23902 27704
rect 23846 24384 23902 24440
rect 25318 55392 25374 55448
rect 24766 54576 24822 54632
rect 24858 53760 24914 53816
rect 25502 52964 25558 53000
rect 25502 52944 25504 52964
rect 25504 52944 25556 52964
rect 25556 52944 25558 52964
rect 25226 52148 25282 52184
rect 25226 52128 25228 52148
rect 25228 52128 25280 52148
rect 25280 52128 25282 52148
rect 25226 51332 25282 51368
rect 25226 51312 25228 51332
rect 25228 51312 25280 51332
rect 25280 51312 25282 51332
rect 25226 50496 25282 50552
rect 25318 49716 25320 49736
rect 25320 49716 25372 49736
rect 25372 49716 25374 49736
rect 23846 19488 23902 19544
rect 23846 17040 23902 17096
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 23294 15408 23350 15464
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23386 13776 23442 13832
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22650 10512 22706 10568
rect 21730 5480 21786 5536
rect 22374 6840 22430 6896
rect 22098 2352 22154 2408
rect 22190 1536 22246 1592
rect 23294 10512 23350 10568
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 23662 6704 23718 6760
rect 23294 5616 23350 5672
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23386 4800 23442 4856
rect 23386 3848 23442 3904
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23294 3476 23296 3496
rect 23296 3476 23348 3496
rect 23348 3476 23350 3496
rect 23294 3440 23350 3476
rect 23386 3168 23442 3224
rect 24858 41384 24914 41440
rect 24766 32544 24822 32600
rect 24490 28464 24546 28520
rect 25318 49680 25374 49716
rect 25226 48864 25282 48920
rect 25226 48084 25228 48104
rect 25228 48084 25280 48104
rect 25280 48084 25282 48104
rect 25226 48048 25282 48084
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 25318 45600 25374 45656
rect 25318 44820 25320 44840
rect 25320 44820 25372 44840
rect 25372 44820 25374 44840
rect 25318 44784 25374 44820
rect 25226 43968 25282 44024
rect 25226 43152 25282 43208
rect 25226 42336 25282 42392
rect 25226 41556 25228 41576
rect 25228 41556 25280 41576
rect 25280 41556 25282 41576
rect 25226 41520 25282 41556
rect 25318 40704 25374 40760
rect 25318 39072 25374 39128
rect 25318 38292 25320 38312
rect 25320 38292 25372 38312
rect 25372 38292 25374 38312
rect 25318 38256 25374 38292
rect 25226 37440 25282 37496
rect 25226 36624 25282 36680
rect 25318 35808 25374 35864
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 25318 34176 25374 34232
rect 25318 33360 25374 33416
rect 25502 39888 25558 39944
rect 24858 29280 24914 29336
rect 24858 26016 24914 26072
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30096 25374 30152
rect 25502 30932 25558 30968
rect 25502 30912 25504 30932
rect 25504 30912 25556 30932
rect 25556 30912 25558 30932
rect 25318 26832 25374 26888
rect 25134 25200 25190 25256
rect 24766 23568 24822 23624
rect 24858 22752 24914 22808
rect 24858 21120 24914 21176
rect 24582 20304 24638 20360
rect 25502 26424 25558 26480
rect 24858 18672 24914 18728
rect 24674 17992 24730 18048
rect 24858 17876 24914 17912
rect 24858 17856 24860 17876
rect 24860 17856 24912 17876
rect 24912 17856 24914 17876
rect 24674 16224 24730 16280
rect 24030 6196 24032 6216
rect 24032 6196 24084 6216
rect 24084 6196 24086 6216
rect 24030 6160 24086 6196
rect 23662 2896 23718 2952
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23938 3984 23994 4040
rect 24858 14592 24914 14648
rect 24766 12960 24822 13016
rect 24858 12144 24914 12200
rect 24858 11328 24914 11384
rect 26330 28056 26386 28112
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 24858 7284 24860 7304
rect 24860 7284 24912 7304
rect 24912 7284 24914 7304
rect 24858 7248 24914 7284
rect 24858 6432 24914 6488
rect 25134 9696 25190 9752
rect 25134 8064 25190 8120
rect 24950 5208 25006 5264
rect 25226 4528 25282 4584
rect 24766 3984 24822 4040
rect 25410 4120 25466 4176
rect 25318 720 25374 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 25313 55450 25379 55453
rect 26200 55450 27000 55480
rect 25313 55448 27000 55450
rect 25313 55392 25318 55448
rect 25374 55392 27000 55448
rect 25313 55390 27000 55392
rect 25313 55387 25379 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 24853 53818 24919 53821
rect 26200 53818 27000 53848
rect 24853 53816 27000 53818
rect 24853 53760 24858 53816
rect 24914 53760 27000 53816
rect 24853 53758 27000 53760
rect 24853 53755 24919 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 25497 53002 25563 53005
rect 26200 53002 27000 53032
rect 25497 53000 27000 53002
rect 25497 52944 25502 53000
rect 25558 52944 27000 53000
rect 25497 52942 27000 52944
rect 25497 52939 25563 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 25221 52186 25287 52189
rect 26200 52186 27000 52216
rect 25221 52184 27000 52186
rect 25221 52128 25226 52184
rect 25282 52128 27000 52184
rect 25221 52126 27000 52128
rect 25221 52123 25287 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25221 51370 25287 51373
rect 26200 51370 27000 51400
rect 25221 51368 27000 51370
rect 25221 51312 25226 51368
rect 25282 51312 27000 51368
rect 25221 51310 27000 51312
rect 25221 51307 25287 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 25221 50554 25287 50557
rect 26200 50554 27000 50584
rect 25221 50552 27000 50554
rect 25221 50496 25226 50552
rect 25282 50496 27000 50552
rect 25221 50494 27000 50496
rect 25221 50491 25287 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49738 25379 49741
rect 26200 49738 27000 49768
rect 25313 49736 27000 49738
rect 25313 49680 25318 49736
rect 25374 49680 27000 49736
rect 25313 49678 27000 49680
rect 25313 49675 25379 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25221 48922 25287 48925
rect 26200 48922 27000 48952
rect 25221 48920 27000 48922
rect 25221 48864 25226 48920
rect 25282 48864 27000 48920
rect 25221 48862 27000 48864
rect 25221 48859 25287 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 25221 48106 25287 48109
rect 26200 48106 27000 48136
rect 25221 48104 27000 48106
rect 25221 48048 25226 48104
rect 25282 48048 27000 48104
rect 25221 48046 27000 48048
rect 25221 48043 25287 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 25221 44026 25287 44029
rect 26200 44026 27000 44056
rect 25221 44024 27000 44026
rect 25221 43968 25226 44024
rect 25282 43968 27000 44024
rect 25221 43966 27000 43968
rect 25221 43963 25287 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 25221 43210 25287 43213
rect 26200 43210 27000 43240
rect 25221 43208 27000 43210
rect 25221 43152 25226 43208
rect 25282 43152 27000 43208
rect 25221 43150 27000 43152
rect 25221 43147 25287 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25221 42394 25287 42397
rect 26200 42394 27000 42424
rect 25221 42392 27000 42394
rect 25221 42336 25226 42392
rect 25282 42336 27000 42392
rect 25221 42334 27000 42336
rect 25221 42331 25287 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25221 41578 25287 41581
rect 26200 41578 27000 41608
rect 25221 41576 27000 41578
rect 25221 41520 25226 41576
rect 25282 41520 27000 41576
rect 25221 41518 27000 41520
rect 25221 41515 25287 41518
rect 26200 41488 27000 41518
rect 23974 41380 23980 41444
rect 24044 41442 24050 41444
rect 24853 41442 24919 41445
rect 24044 41440 24919 41442
rect 24044 41384 24858 41440
rect 24914 41384 24919 41440
rect 24044 41382 24919 41384
rect 24044 41380 24050 41382
rect 24853 41379 24919 41382
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 25497 39946 25563 39949
rect 26200 39946 27000 39976
rect 25497 39944 27000 39946
rect 25497 39888 25502 39944
rect 25558 39888 27000 39944
rect 25497 39886 27000 39888
rect 25497 39883 25563 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25221 37498 25287 37501
rect 26200 37498 27000 37528
rect 25221 37496 27000 37498
rect 25221 37440 25226 37496
rect 25282 37440 27000 37496
rect 25221 37438 27000 37440
rect 25221 37435 25287 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 25221 36682 25287 36685
rect 26200 36682 27000 36712
rect 25221 36680 27000 36682
rect 25221 36624 25226 36680
rect 25282 36624 27000 36680
rect 25221 36622 27000 36624
rect 25221 36619 25287 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 21081 35594 21147 35597
rect 22134 35594 22140 35596
rect 21081 35592 22140 35594
rect 21081 35536 21086 35592
rect 21142 35536 22140 35592
rect 21081 35534 22140 35536
rect 21081 35531 21147 35534
rect 22134 35532 22140 35534
rect 22204 35532 22210 35596
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 25313 33418 25379 33421
rect 26200 33418 27000 33448
rect 25313 33416 27000 33418
rect 25313 33360 25318 33416
rect 25374 33360 27000 33416
rect 25313 33358 27000 33360
rect 25313 33355 25379 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 22134 33084 22140 33148
rect 22204 33146 22210 33148
rect 22645 33146 22711 33149
rect 22204 33144 22711 33146
rect 22204 33088 22650 33144
rect 22706 33088 22711 33144
rect 22204 33086 22711 33088
rect 22204 33084 22210 33086
rect 22645 33083 22711 33086
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 24761 32602 24827 32605
rect 26200 32602 27000 32632
rect 24761 32600 27000 32602
rect 24761 32544 24766 32600
rect 24822 32544 27000 32600
rect 24761 32542 27000 32544
rect 24761 32539 24827 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25497 30970 25563 30973
rect 26200 30970 27000 31000
rect 25497 30968 27000 30970
rect 25497 30912 25502 30968
rect 25558 30912 27000 30968
rect 25497 30910 27000 30912
rect 25497 30907 25563 30910
rect 26200 30880 27000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 24853 29338 24919 29341
rect 26200 29338 27000 29368
rect 24853 29336 27000 29338
rect 24853 29280 24858 29336
rect 24914 29280 27000 29336
rect 24853 29278 27000 29280
rect 24853 29275 24919 29278
rect 26200 29248 27000 29278
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24485 28522 24551 28525
rect 26200 28522 27000 28552
rect 24485 28520 27000 28522
rect 24485 28464 24490 28520
rect 24546 28464 27000 28520
rect 24485 28462 27000 28464
rect 24485 28459 24551 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 16113 28114 16179 28117
rect 26325 28114 26391 28117
rect 16113 28112 26391 28114
rect 16113 28056 16118 28112
rect 16174 28056 26330 28112
rect 26386 28056 26391 28112
rect 16113 28054 26391 28056
rect 16113 28051 16179 28054
rect 26325 28051 26391 28054
rect 18505 27844 18571 27845
rect 18454 27780 18460 27844
rect 18524 27842 18571 27844
rect 18524 27840 18616 27842
rect 18566 27784 18616 27840
rect 18524 27782 18616 27784
rect 18524 27780 18571 27782
rect 18505 27779 18571 27780
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 23841 27706 23907 27709
rect 26200 27706 27000 27736
rect 23841 27704 27000 27706
rect 23841 27648 23846 27704
rect 23902 27648 27000 27704
rect 23841 27646 27000 27648
rect 23841 27643 23907 27646
rect 26200 27616 27000 27646
rect 15561 27298 15627 27301
rect 15694 27298 15700 27300
rect 15561 27296 15700 27298
rect 15561 27240 15566 27296
rect 15622 27240 15700 27296
rect 15561 27238 15700 27240
rect 15561 27235 15627 27238
rect 15694 27236 15700 27238
rect 15764 27236 15770 27300
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25313 26890 25379 26893
rect 26200 26890 27000 26920
rect 25313 26888 27000 26890
rect 25313 26832 25318 26888
rect 25374 26832 27000 26888
rect 25313 26830 27000 26832
rect 25313 26827 25379 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 20345 26482 20411 26485
rect 25497 26482 25563 26485
rect 20345 26480 25563 26482
rect 20345 26424 20350 26480
rect 20406 26424 25502 26480
rect 25558 26424 25563 26480
rect 20345 26422 25563 26424
rect 20345 26419 20411 26422
rect 25497 26419 25563 26422
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 24853 26074 24919 26077
rect 26200 26074 27000 26104
rect 24853 26072 27000 26074
rect 24853 26016 24858 26072
rect 24914 26016 27000 26072
rect 24853 26014 27000 26016
rect 24853 26011 24919 26014
rect 26200 25984 27000 26014
rect 17401 25802 17467 25805
rect 17718 25802 17724 25804
rect 17401 25800 17724 25802
rect 17401 25744 17406 25800
rect 17462 25744 17724 25800
rect 17401 25742 17724 25744
rect 17401 25739 17467 25742
rect 17718 25740 17724 25742
rect 17788 25740 17794 25804
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 19374 24924 19380 24988
rect 19444 24986 19450 24988
rect 19701 24986 19767 24989
rect 19444 24984 19767 24986
rect 19444 24928 19706 24984
rect 19762 24928 19767 24984
rect 19444 24926 19767 24928
rect 19444 24924 19450 24926
rect 19701 24923 19767 24926
rect 15193 24714 15259 24717
rect 16430 24714 16436 24716
rect 15193 24712 16436 24714
rect 15193 24656 15198 24712
rect 15254 24656 16436 24712
rect 15193 24654 16436 24656
rect 15193 24651 15259 24654
rect 16430 24652 16436 24654
rect 16500 24652 16506 24716
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 23841 24442 23907 24445
rect 26200 24442 27000 24472
rect 23841 24440 27000 24442
rect 23841 24384 23846 24440
rect 23902 24384 27000 24440
rect 23841 24382 27000 24384
rect 23841 24379 23907 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 24761 23626 24827 23629
rect 26200 23626 27000 23656
rect 24761 23624 27000 23626
rect 24761 23568 24766 23624
rect 24822 23568 27000 23624
rect 24761 23566 27000 23568
rect 24761 23563 24827 23566
rect 26200 23536 27000 23566
rect 19057 23490 19123 23493
rect 19977 23490 20043 23493
rect 19057 23488 20043 23490
rect 19057 23432 19062 23488
rect 19118 23432 19982 23488
rect 20038 23432 20043 23488
rect 19057 23430 20043 23432
rect 19057 23427 19123 23430
rect 19977 23427 20043 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 17309 22812 17375 22813
rect 17309 22808 17356 22812
rect 17420 22810 17426 22812
rect 24853 22810 24919 22813
rect 26200 22810 27000 22840
rect 17309 22752 17314 22808
rect 17309 22748 17356 22752
rect 17420 22750 17466 22810
rect 24853 22808 27000 22810
rect 24853 22752 24858 22808
rect 24914 22752 27000 22808
rect 24853 22750 27000 22752
rect 17420 22748 17426 22750
rect 17309 22747 17375 22748
rect 24853 22747 24919 22750
rect 26200 22720 27000 22750
rect 20437 22404 20503 22405
rect 20437 22402 20484 22404
rect 20392 22400 20484 22402
rect 20392 22344 20442 22400
rect 20392 22342 20484 22344
rect 20437 22340 20484 22342
rect 20548 22340 20554 22404
rect 20437 22339 20503 22340
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 19057 22266 19123 22269
rect 18830 22264 19123 22266
rect 18830 22208 19062 22264
rect 19118 22208 19123 22264
rect 18830 22206 19123 22208
rect 18689 22130 18755 22133
rect 18830 22130 18890 22206
rect 19057 22203 19123 22206
rect 18689 22128 18890 22130
rect 18689 22072 18694 22128
rect 18750 22072 18890 22128
rect 18689 22070 18890 22072
rect 18689 22067 18755 22070
rect 22829 21994 22895 21997
rect 26200 21994 27000 22024
rect 22829 21992 27000 21994
rect 22829 21936 22834 21992
rect 22890 21936 27000 21992
rect 22829 21934 27000 21936
rect 22829 21931 22895 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 24853 21178 24919 21181
rect 26200 21178 27000 21208
rect 24853 21176 27000 21178
rect 24853 21120 24858 21176
rect 24914 21120 27000 21176
rect 24853 21118 27000 21120
rect 24853 21115 24919 21118
rect 26200 21088 27000 21118
rect 13670 20844 13676 20908
rect 13740 20906 13746 20908
rect 19374 20906 19380 20908
rect 13740 20846 19380 20906
rect 13740 20844 13746 20846
rect 19374 20844 19380 20846
rect 19444 20844 19450 20908
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 24577 20362 24643 20365
rect 26200 20362 27000 20392
rect 24577 20360 27000 20362
rect 24577 20304 24582 20360
rect 24638 20304 27000 20360
rect 24577 20302 27000 20304
rect 24577 20299 24643 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 23841 19546 23907 19549
rect 26200 19546 27000 19576
rect 23841 19544 27000 19546
rect 23841 19488 23846 19544
rect 23902 19488 27000 19544
rect 23841 19486 27000 19488
rect 23841 19483 23907 19486
rect 26200 19456 27000 19486
rect 19558 19348 19564 19412
rect 19628 19410 19634 19412
rect 19701 19410 19767 19413
rect 19628 19408 19767 19410
rect 19628 19352 19706 19408
rect 19762 19352 19767 19408
rect 19628 19350 19767 19352
rect 19628 19348 19634 19350
rect 19701 19347 19767 19350
rect 18965 19274 19031 19277
rect 23422 19274 23428 19276
rect 18965 19272 23428 19274
rect 18965 19216 18970 19272
rect 19026 19216 23428 19272
rect 18965 19214 23428 19216
rect 18965 19211 19031 19214
rect 23422 19212 23428 19214
rect 23492 19212 23498 19276
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 24853 18730 24919 18733
rect 26200 18730 27000 18760
rect 24853 18728 27000 18730
rect 24853 18672 24858 18728
rect 24914 18672 27000 18728
rect 24853 18670 27000 18672
rect 24853 18667 24919 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 21081 18050 21147 18053
rect 24669 18052 24735 18053
rect 21214 18050 21220 18052
rect 21081 18048 21220 18050
rect 21081 17992 21086 18048
rect 21142 17992 21220 18048
rect 21081 17990 21220 17992
rect 21081 17987 21147 17990
rect 21214 17988 21220 17990
rect 21284 17988 21290 18052
rect 24669 18048 24716 18052
rect 24780 18050 24786 18052
rect 24669 17992 24674 18048
rect 24669 17988 24716 17992
rect 24780 17990 24826 18050
rect 24780 17988 24786 17990
rect 24669 17987 24735 17988
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 17718 17852 17724 17916
rect 17788 17914 17794 17916
rect 17861 17914 17927 17917
rect 17788 17912 17927 17914
rect 17788 17856 17866 17912
rect 17922 17856 17927 17912
rect 17788 17854 17927 17856
rect 17788 17852 17794 17854
rect 17861 17851 17927 17854
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 23841 17098 23907 17101
rect 26200 17098 27000 17128
rect 23841 17096 27000 17098
rect 23841 17040 23846 17096
rect 23902 17040 27000 17096
rect 23841 17038 27000 17040
rect 23841 17035 23907 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 21766 16628 21772 16692
rect 21836 16690 21842 16692
rect 21909 16690 21975 16693
rect 21836 16688 21975 16690
rect 21836 16632 21914 16688
rect 21970 16632 21975 16688
rect 21836 16630 21975 16632
rect 21836 16628 21842 16630
rect 21909 16627 21975 16630
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 17309 16284 17375 16285
rect 17309 16282 17356 16284
rect 17264 16280 17356 16282
rect 17264 16224 17314 16280
rect 17264 16222 17356 16224
rect 17309 16220 17356 16222
rect 17420 16220 17426 16284
rect 24669 16282 24735 16285
rect 26200 16282 27000 16312
rect 24669 16280 27000 16282
rect 24669 16224 24674 16280
rect 24730 16224 27000 16280
rect 24669 16222 27000 16224
rect 17309 16219 17375 16220
rect 24669 16219 24735 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 23289 15466 23355 15469
rect 26200 15466 27000 15496
rect 23289 15464 27000 15466
rect 23289 15408 23294 15464
rect 23350 15408 27000 15464
rect 23289 15406 27000 15408
rect 23289 15403 23355 15406
rect 26200 15376 27000 15406
rect 17217 15330 17283 15333
rect 17350 15330 17356 15332
rect 17217 15328 17356 15330
rect 17217 15272 17222 15328
rect 17278 15272 17356 15328
rect 17217 15270 17356 15272
rect 17217 15267 17283 15270
rect 17350 15268 17356 15270
rect 17420 15268 17426 15332
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24853 14650 24919 14653
rect 26200 14650 27000 14680
rect 24853 14648 27000 14650
rect 24853 14592 24858 14648
rect 24914 14592 27000 14648
rect 24853 14590 27000 14592
rect 24853 14587 24919 14590
rect 26200 14560 27000 14590
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 12566 13908 12572 13972
rect 12636 13970 12642 13972
rect 13813 13970 13879 13973
rect 12636 13968 13879 13970
rect 12636 13912 13818 13968
rect 13874 13912 13879 13968
rect 12636 13910 13879 13912
rect 12636 13908 12642 13910
rect 13813 13907 13879 13910
rect 23381 13834 23447 13837
rect 26200 13834 27000 13864
rect 23381 13832 27000 13834
rect 23381 13776 23386 13832
rect 23442 13776 27000 13832
rect 23381 13774 27000 13776
rect 23381 13771 23447 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 24761 13018 24827 13021
rect 26200 13018 27000 13048
rect 24761 13016 27000 13018
rect 24761 12960 24766 13016
rect 24822 12960 27000 13016
rect 24761 12958 27000 12960
rect 24761 12955 24827 12958
rect 26200 12928 27000 12958
rect 15377 12610 15443 12613
rect 15745 12610 15811 12613
rect 15377 12608 15811 12610
rect 15377 12552 15382 12608
rect 15438 12552 15750 12608
rect 15806 12552 15811 12608
rect 15377 12550 15811 12552
rect 15377 12547 15443 12550
rect 15745 12547 15811 12550
rect 16798 12548 16804 12612
rect 16868 12610 16874 12612
rect 17217 12610 17283 12613
rect 16868 12608 17283 12610
rect 16868 12552 17222 12608
rect 17278 12552 17283 12608
rect 16868 12550 17283 12552
rect 16868 12548 16874 12550
rect 17217 12547 17283 12550
rect 18413 12610 18479 12613
rect 18781 12610 18847 12613
rect 18413 12608 18847 12610
rect 18413 12552 18418 12608
rect 18474 12552 18786 12608
rect 18842 12552 18847 12608
rect 18413 12550 18847 12552
rect 18413 12547 18479 12550
rect 18781 12547 18847 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 12433 12474 12499 12477
rect 12709 12474 12775 12477
rect 12433 12472 12775 12474
rect 12433 12416 12438 12472
rect 12494 12416 12714 12472
rect 12770 12416 12775 12472
rect 12433 12414 12775 12416
rect 12433 12411 12499 12414
rect 12709 12411 12775 12414
rect 14273 12474 14339 12477
rect 14733 12474 14799 12477
rect 14273 12472 14799 12474
rect 14273 12416 14278 12472
rect 14334 12416 14738 12472
rect 14794 12416 14799 12472
rect 14273 12414 14799 12416
rect 14273 12411 14339 12414
rect 14733 12411 14799 12414
rect 24853 12202 24919 12205
rect 26200 12202 27000 12232
rect 24853 12200 27000 12202
rect 24853 12144 24858 12200
rect 24914 12144 27000 12200
rect 24853 12142 27000 12144
rect 24853 12139 24919 12142
rect 26200 12112 27000 12142
rect 21449 12066 21515 12069
rect 23974 12066 23980 12068
rect 21449 12064 23980 12066
rect 21449 12008 21454 12064
rect 21510 12008 23980 12064
rect 21449 12006 23980 12008
rect 21449 12003 21515 12006
rect 23974 12004 23980 12006
rect 24044 12004 24050 12068
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 12065 11658 12131 11661
rect 13077 11658 13143 11661
rect 12065 11656 13143 11658
rect 12065 11600 12070 11656
rect 12126 11600 13082 11656
rect 13138 11600 13143 11656
rect 12065 11598 13143 11600
rect 12065 11595 12131 11598
rect 13077 11595 13143 11598
rect 14641 11524 14707 11525
rect 14590 11522 14596 11524
rect 14550 11462 14596 11522
rect 14660 11520 14707 11524
rect 14702 11464 14707 11520
rect 14590 11460 14596 11462
rect 14660 11460 14707 11464
rect 14641 11459 14707 11460
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 17677 10706 17743 10709
rect 19558 10706 19564 10708
rect 17677 10704 19564 10706
rect 17677 10648 17682 10704
rect 17738 10648 19564 10704
rect 17677 10646 19564 10648
rect 17677 10643 17743 10646
rect 19558 10644 19564 10646
rect 19628 10644 19634 10708
rect 17677 10570 17743 10573
rect 18965 10570 19031 10573
rect 17677 10568 19031 10570
rect 17677 10512 17682 10568
rect 17738 10512 18970 10568
rect 19026 10512 19031 10568
rect 17677 10510 19031 10512
rect 17677 10507 17743 10510
rect 18965 10507 19031 10510
rect 19609 10570 19675 10573
rect 22645 10570 22711 10573
rect 19609 10568 22711 10570
rect 19609 10512 19614 10568
rect 19670 10512 22650 10568
rect 22706 10512 22711 10568
rect 19609 10510 22711 10512
rect 19609 10507 19675 10510
rect 22645 10507 22711 10510
rect 23289 10570 23355 10573
rect 26200 10570 27000 10600
rect 23289 10568 27000 10570
rect 23289 10512 23294 10568
rect 23350 10512 27000 10568
rect 23289 10510 27000 10512
rect 23289 10507 23355 10510
rect 26200 10480 27000 10510
rect 14089 10436 14155 10437
rect 14038 10434 14044 10436
rect 13962 10374 14044 10434
rect 14108 10434 14155 10436
rect 15694 10434 15700 10436
rect 14108 10432 15700 10434
rect 14150 10376 15700 10432
rect 14038 10372 14044 10374
rect 14108 10374 15700 10376
rect 14108 10372 14155 10374
rect 15694 10372 15700 10374
rect 15764 10434 15770 10436
rect 20437 10434 20503 10437
rect 22461 10434 22527 10437
rect 15764 10432 22527 10434
rect 15764 10376 20442 10432
rect 20498 10376 22466 10432
rect 22522 10376 22527 10432
rect 15764 10374 22527 10376
rect 15764 10372 15770 10374
rect 14089 10371 14155 10372
rect 20437 10371 20503 10374
rect 22461 10371 22527 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 18413 10164 18479 10165
rect 18413 10162 18460 10164
rect 18368 10160 18460 10162
rect 18368 10104 18418 10160
rect 18368 10102 18460 10104
rect 18413 10100 18460 10102
rect 18524 10100 18530 10164
rect 18413 10099 18479 10100
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 25129 9754 25195 9757
rect 26200 9754 27000 9784
rect 25129 9752 27000 9754
rect 25129 9696 25134 9752
rect 25190 9696 27000 9752
rect 25129 9694 27000 9696
rect 25129 9691 25195 9694
rect 26200 9664 27000 9694
rect 19149 9618 19215 9621
rect 21214 9618 21220 9620
rect 19149 9616 21220 9618
rect 19149 9560 19154 9616
rect 19210 9560 21220 9616
rect 19149 9558 21220 9560
rect 19149 9555 19215 9558
rect 21214 9556 21220 9558
rect 21284 9556 21290 9620
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 5349 9210 5415 9213
rect 12382 9210 12388 9212
rect 5349 9208 12388 9210
rect 5349 9152 5354 9208
rect 5410 9152 12388 9208
rect 5349 9150 12388 9152
rect 5349 9147 5415 9150
rect 12382 9148 12388 9150
rect 12452 9148 12458 9212
rect 13537 8938 13603 8941
rect 17033 8938 17099 8941
rect 13537 8936 17099 8938
rect 13537 8880 13542 8936
rect 13598 8880 17038 8936
rect 17094 8880 17099 8936
rect 13537 8878 17099 8880
rect 13537 8875 13603 8878
rect 17033 8875 17099 8878
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 0 8802 800 8832
rect 3877 8802 3943 8805
rect 0 8800 3943 8802
rect 0 8744 3882 8800
rect 3938 8744 3943 8800
rect 0 8742 3943 8744
rect 0 8712 800 8742
rect 3877 8739 3943 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 12801 8530 12867 8533
rect 17309 8530 17375 8533
rect 12801 8528 17375 8530
rect 12801 8472 12806 8528
rect 12862 8472 17314 8528
rect 17370 8472 17375 8528
rect 12801 8470 17375 8472
rect 12801 8467 12867 8470
rect 17309 8467 17375 8470
rect 14406 8332 14412 8396
rect 14476 8394 14482 8396
rect 16205 8394 16271 8397
rect 14476 8392 16271 8394
rect 14476 8336 16210 8392
rect 16266 8336 16271 8392
rect 14476 8334 16271 8336
rect 14476 8332 14482 8334
rect 16205 8331 16271 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 11789 7986 11855 7989
rect 16798 7986 16804 7988
rect 11789 7984 16804 7986
rect 11789 7928 11794 7984
rect 11850 7928 16804 7984
rect 11789 7926 16804 7928
rect 11789 7923 11855 7926
rect 16798 7924 16804 7926
rect 16868 7924 16874 7988
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 14365 6898 14431 6901
rect 14590 6898 14596 6900
rect 14365 6896 14596 6898
rect 14365 6840 14370 6896
rect 14426 6840 14596 6896
rect 14365 6838 14596 6840
rect 14365 6835 14431 6838
rect 14590 6836 14596 6838
rect 14660 6836 14666 6900
rect 17309 6898 17375 6901
rect 22369 6898 22435 6901
rect 17309 6896 22435 6898
rect 17309 6840 17314 6896
rect 17370 6840 22374 6896
rect 22430 6840 22435 6896
rect 17309 6838 22435 6840
rect 17309 6835 17375 6838
rect 22369 6835 22435 6838
rect 13629 6762 13695 6765
rect 23657 6762 23723 6765
rect 13629 6760 23723 6762
rect 13629 6704 13634 6760
rect 13690 6704 23662 6760
rect 23718 6704 23723 6760
rect 13629 6702 23723 6704
rect 13629 6699 13695 6702
rect 23657 6699 23723 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 4061 6490 4127 6493
rect 14089 6492 14155 6493
rect 0 6488 4127 6490
rect 0 6432 4066 6488
rect 4122 6432 4127 6488
rect 0 6430 4127 6432
rect 0 6400 800 6430
rect 4061 6427 4127 6430
rect 14038 6428 14044 6492
rect 14108 6490 14155 6492
rect 24853 6490 24919 6493
rect 26200 6490 27000 6520
rect 14108 6488 14200 6490
rect 14150 6432 14200 6488
rect 14108 6430 14200 6432
rect 24853 6488 27000 6490
rect 24853 6432 24858 6488
rect 24914 6432 27000 6488
rect 24853 6430 27000 6432
rect 14108 6428 14155 6430
rect 14089 6427 14155 6428
rect 24853 6427 24919 6430
rect 26200 6400 27000 6430
rect 10225 6218 10291 6221
rect 24025 6218 24091 6221
rect 10225 6216 24091 6218
rect 10225 6160 10230 6216
rect 10286 6160 24030 6216
rect 24086 6160 24091 6216
rect 10225 6158 24091 6160
rect 10225 6155 10291 6158
rect 24025 6155 24091 6158
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 12249 5810 12315 5813
rect 17309 5810 17375 5813
rect 12249 5808 17375 5810
rect 12249 5752 12254 5808
rect 12310 5752 17314 5808
rect 17370 5752 17375 5808
rect 12249 5750 17375 5752
rect 12249 5747 12315 5750
rect 17309 5747 17375 5750
rect 15285 5674 15351 5677
rect 16430 5674 16436 5676
rect 15285 5672 16436 5674
rect 15285 5616 15290 5672
rect 15346 5616 16436 5672
rect 15285 5614 16436 5616
rect 15285 5611 15351 5614
rect 16430 5612 16436 5614
rect 16500 5674 16506 5676
rect 20069 5674 20135 5677
rect 21265 5674 21331 5677
rect 16500 5672 21331 5674
rect 16500 5616 20074 5672
rect 20130 5616 21270 5672
rect 21326 5616 21331 5672
rect 16500 5614 21331 5616
rect 16500 5612 16506 5614
rect 20069 5611 20135 5614
rect 21265 5611 21331 5614
rect 23289 5674 23355 5677
rect 26200 5674 27000 5704
rect 23289 5672 27000 5674
rect 23289 5616 23294 5672
rect 23350 5616 27000 5672
rect 23289 5614 27000 5616
rect 23289 5611 23355 5614
rect 26200 5584 27000 5614
rect 21725 5540 21791 5541
rect 21725 5536 21772 5540
rect 21836 5538 21842 5540
rect 21725 5480 21730 5536
rect 21725 5476 21772 5480
rect 21836 5478 21882 5538
rect 21836 5476 21842 5478
rect 21725 5475 21791 5476
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 12249 5402 12315 5405
rect 17677 5402 17743 5405
rect 12249 5400 17743 5402
rect 12249 5344 12254 5400
rect 12310 5344 17682 5400
rect 17738 5344 17743 5400
rect 12249 5342 17743 5344
rect 12249 5339 12315 5342
rect 17677 5339 17743 5342
rect 12893 5266 12959 5269
rect 24945 5266 25011 5269
rect 12893 5264 25011 5266
rect 12893 5208 12898 5264
rect 12954 5208 24950 5264
rect 25006 5208 25011 5264
rect 12893 5206 25011 5208
rect 12893 5203 12959 5206
rect 24945 5203 25011 5206
rect 11145 5130 11211 5133
rect 20897 5130 20963 5133
rect 11145 5128 20963 5130
rect 11145 5072 11150 5128
rect 11206 5072 20902 5128
rect 20958 5072 20963 5128
rect 11145 5070 20963 5072
rect 11145 5067 11211 5070
rect 20897 5067 20963 5070
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 11145 4586 11211 4589
rect 25221 4586 25287 4589
rect 11145 4584 25287 4586
rect 11145 4528 11150 4584
rect 11206 4528 25226 4584
rect 25282 4528 25287 4584
rect 11145 4526 25287 4528
rect 11145 4523 11211 4526
rect 25221 4523 25287 4526
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4178 800 4208
rect 25405 4178 25471 4181
rect 0 4176 25471 4178
rect 0 4120 25410 4176
rect 25466 4120 25471 4176
rect 0 4118 25471 4120
rect 0 4088 800 4118
rect 25405 4115 25471 4118
rect 5165 4042 5231 4045
rect 11237 4042 11303 4045
rect 5165 4040 11303 4042
rect 5165 3984 5170 4040
rect 5226 3984 11242 4040
rect 11298 3984 11303 4040
rect 5165 3982 11303 3984
rect 5165 3979 5231 3982
rect 11237 3979 11303 3982
rect 12801 4042 12867 4045
rect 14365 4044 14431 4045
rect 13670 4042 13676 4044
rect 12801 4040 13676 4042
rect 12801 3984 12806 4040
rect 12862 3984 13676 4040
rect 12801 3982 13676 3984
rect 12801 3979 12867 3982
rect 13670 3980 13676 3982
rect 13740 3980 13746 4044
rect 14365 4042 14412 4044
rect 14320 4040 14412 4042
rect 14320 3984 14370 4040
rect 14320 3982 14412 3984
rect 14365 3980 14412 3982
rect 14476 3980 14482 4044
rect 23422 3980 23428 4044
rect 23492 4042 23498 4044
rect 23933 4042 23999 4045
rect 24761 4044 24827 4045
rect 23492 4040 23999 4042
rect 23492 3984 23938 4040
rect 23994 3984 23999 4040
rect 23492 3982 23999 3984
rect 23492 3980 23498 3982
rect 14365 3979 14431 3980
rect 23933 3979 23999 3982
rect 24710 3980 24716 4044
rect 24780 4042 24827 4044
rect 26200 4042 27000 4072
rect 24780 4040 24872 4042
rect 24822 3984 24872 4040
rect 24780 3982 24872 3984
rect 25086 3982 27000 4042
rect 24780 3980 24827 3982
rect 24761 3979 24827 3980
rect 23381 3906 23447 3909
rect 25086 3906 25146 3982
rect 26200 3952 27000 3982
rect 23381 3904 25146 3906
rect 23381 3848 23386 3904
rect 23442 3848 25146 3904
rect 23381 3846 25146 3848
rect 23381 3843 23447 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 15653 3634 15719 3637
rect 17350 3634 17356 3636
rect 15653 3632 17356 3634
rect 15653 3576 15658 3632
rect 15714 3576 17356 3632
rect 15653 3574 17356 3576
rect 15653 3571 15719 3574
rect 17350 3572 17356 3574
rect 17420 3572 17426 3636
rect 7925 3498 7991 3501
rect 23289 3498 23355 3501
rect 7925 3496 23355 3498
rect 7925 3440 7930 3496
rect 7986 3440 23294 3496
rect 23350 3440 23355 3496
rect 7925 3438 23355 3440
rect 7925 3435 7991 3438
rect 23289 3435 23355 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 23381 3226 23447 3229
rect 26200 3226 27000 3256
rect 23381 3224 27000 3226
rect 23381 3168 23386 3224
rect 23442 3168 27000 3224
rect 23381 3166 27000 3168
rect 23381 3163 23447 3166
rect 26200 3136 27000 3166
rect 5717 3090 5783 3093
rect 13353 3090 13419 3093
rect 5717 3088 13419 3090
rect 5717 3032 5722 3088
rect 5778 3032 13358 3088
rect 13414 3032 13419 3088
rect 5717 3030 13419 3032
rect 5717 3027 5783 3030
rect 13353 3027 13419 3030
rect 13445 2954 13511 2957
rect 23657 2954 23723 2957
rect 13445 2952 23723 2954
rect 13445 2896 13450 2952
rect 13506 2896 23662 2952
rect 23718 2896 23723 2952
rect 13445 2894 23723 2896
rect 13445 2891 13511 2894
rect 23657 2891 23723 2894
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 22093 2410 22159 2413
rect 26200 2410 27000 2440
rect 22093 2408 27000 2410
rect 22093 2352 22098 2408
rect 22154 2352 27000 2408
rect 22093 2350 27000 2352
rect 22093 2347 22159 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 20478 1866 20484 1868
rect 0 1806 20484 1866
rect 0 1776 800 1806
rect 20478 1804 20484 1806
rect 20548 1804 20554 1868
rect 22185 1594 22251 1597
rect 26200 1594 27000 1624
rect 22185 1592 27000 1594
rect 22185 1536 22190 1592
rect 22246 1536 27000 1592
rect 22185 1534 27000 1536
rect 22185 1531 22251 1534
rect 26200 1504 27000 1534
rect 25313 778 25379 781
rect 26200 778 27000 808
rect 25313 776 27000 778
rect 25313 720 25318 776
rect 25374 720 27000 776
rect 25313 718 27000 720
rect 25313 715 25379 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 23980 41380 24044 41444
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 22140 35532 22204 35596
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 22140 33084 22204 33148
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 18460 27840 18524 27844
rect 18460 27784 18510 27840
rect 18510 27784 18524 27840
rect 18460 27780 18524 27784
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 15700 27236 15764 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 17724 25740 17788 25804
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 19380 24924 19444 24988
rect 16436 24652 16500 24716
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 17356 22808 17420 22812
rect 17356 22752 17370 22808
rect 17370 22752 17420 22808
rect 17356 22748 17420 22752
rect 20484 22400 20548 22404
rect 20484 22344 20498 22400
rect 20498 22344 20548 22400
rect 20484 22340 20548 22344
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 13676 20844 13740 20908
rect 19380 20844 19444 20908
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 19564 19348 19628 19412
rect 23428 19212 23492 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 21220 17988 21284 18052
rect 24716 18048 24780 18052
rect 24716 17992 24730 18048
rect 24730 17992 24780 18048
rect 24716 17988 24780 17992
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 17724 17852 17788 17916
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 21772 16628 21836 16692
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 17356 16280 17420 16284
rect 17356 16224 17370 16280
rect 17370 16224 17420 16280
rect 17356 16220 17420 16224
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 17356 15268 17420 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 12572 13908 12636 13972
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 16804 12548 16868 12612
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 23980 12004 24044 12068
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 14596 11520 14660 11524
rect 14596 11464 14646 11520
rect 14646 11464 14660 11520
rect 14596 11460 14660 11464
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 19564 10644 19628 10708
rect 14044 10432 14108 10436
rect 14044 10376 14094 10432
rect 14094 10376 14108 10432
rect 14044 10372 14108 10376
rect 15700 10372 15764 10436
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 18460 10160 18524 10164
rect 18460 10104 18474 10160
rect 18474 10104 18524 10160
rect 18460 10100 18524 10104
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 21220 9556 21284 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 12388 9148 12452 9212
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 14412 8332 14476 8396
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 16804 7924 16868 7988
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 14596 6836 14660 6900
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 14044 6488 14108 6492
rect 14044 6432 14094 6488
rect 14094 6432 14108 6488
rect 14044 6428 14108 6432
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 16436 5612 16500 5676
rect 21772 5536 21836 5540
rect 21772 5480 21786 5536
rect 21786 5480 21836 5536
rect 21772 5476 21836 5480
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 13676 3980 13740 4044
rect 14412 4040 14476 4044
rect 14412 3984 14426 4040
rect 14426 3984 14476 4040
rect 14412 3980 14476 3984
rect 23428 3980 23492 4044
rect 24716 4040 24780 4044
rect 24716 3984 24766 4040
rect 24766 3984 24780 4040
rect 24716 3980 24780 3984
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 17356 3572 17420 3636
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 20484 1804 20548 1868
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 23979 41444 24045 41445
rect 23979 41380 23980 41444
rect 24044 41380 24045 41444
rect 23979 41379 24045 41380
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22139 35596 22205 35597
rect 22139 35532 22140 35596
rect 22204 35532 22205 35596
rect 22139 35531 22205 35532
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 22142 33149 22202 35531
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22139 33148 22205 33149
rect 22139 33084 22140 33148
rect 22204 33084 22205 33148
rect 22139 33083 22205 33084
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 15699 27300 15765 27301
rect 15699 27236 15700 27300
rect 15764 27236 15765 27300
rect 15699 27235 15765 27236
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 13675 20908 13741 20909
rect 13675 20844 13676 20908
rect 13740 20844 13741 20908
rect 13675 20843 13741 20844
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12571 13972 12637 13973
rect 12571 13908 12572 13972
rect 12636 13908 12637 13972
rect 12571 13907 12637 13908
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 12387 9212 12453 9213
rect 12387 9148 12388 9212
rect 12452 9210 12453 9212
rect 12574 9210 12634 13907
rect 12452 9150 12634 9210
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12452 9148 12453 9150
rect 12387 9147 12453 9148
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 13678 4045 13738 20843
rect 14595 11524 14661 11525
rect 14595 11460 14596 11524
rect 14660 11460 14661 11524
rect 14595 11459 14661 11460
rect 14043 10436 14109 10437
rect 14043 10372 14044 10436
rect 14108 10372 14109 10436
rect 14043 10371 14109 10372
rect 14046 6493 14106 10371
rect 14411 8396 14477 8397
rect 14411 8332 14412 8396
rect 14476 8332 14477 8396
rect 14411 8331 14477 8332
rect 14043 6492 14109 6493
rect 14043 6428 14044 6492
rect 14108 6428 14109 6492
rect 14043 6427 14109 6428
rect 14414 4045 14474 8331
rect 14598 6901 14658 11459
rect 15702 10437 15762 27235
rect 17944 27232 18264 28256
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 18459 27844 18525 27845
rect 18459 27780 18460 27844
rect 18524 27780 18525 27844
rect 18459 27779 18525 27780
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17723 25804 17789 25805
rect 17723 25740 17724 25804
rect 17788 25740 17789 25804
rect 17723 25739 17789 25740
rect 16435 24716 16501 24717
rect 16435 24652 16436 24716
rect 16500 24652 16501 24716
rect 16435 24651 16501 24652
rect 15699 10436 15765 10437
rect 15699 10372 15700 10436
rect 15764 10372 15765 10436
rect 15699 10371 15765 10372
rect 14595 6900 14661 6901
rect 14595 6836 14596 6900
rect 14660 6836 14661 6900
rect 14595 6835 14661 6836
rect 16438 5677 16498 24651
rect 17355 22812 17421 22813
rect 17355 22748 17356 22812
rect 17420 22748 17421 22812
rect 17355 22747 17421 22748
rect 17358 16285 17418 22747
rect 17726 17917 17786 25739
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17723 17916 17789 17917
rect 17723 17852 17724 17916
rect 17788 17852 17789 17916
rect 17723 17851 17789 17852
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17355 16284 17421 16285
rect 17355 16220 17356 16284
rect 17420 16220 17421 16284
rect 17355 16219 17421 16220
rect 17355 15332 17421 15333
rect 17355 15268 17356 15332
rect 17420 15268 17421 15332
rect 17355 15267 17421 15268
rect 16803 12612 16869 12613
rect 16803 12548 16804 12612
rect 16868 12548 16869 12612
rect 16803 12547 16869 12548
rect 16806 7989 16866 12547
rect 16803 7988 16869 7989
rect 16803 7924 16804 7988
rect 16868 7924 16869 7988
rect 16803 7923 16869 7924
rect 16435 5676 16501 5677
rect 16435 5612 16436 5676
rect 16500 5612 16501 5676
rect 16435 5611 16501 5612
rect 13675 4044 13741 4045
rect 13675 3980 13676 4044
rect 13740 3980 13741 4044
rect 13675 3979 13741 3980
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 17358 3637 17418 15267
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 18462 10165 18522 27779
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 19379 24988 19445 24989
rect 19379 24924 19380 24988
rect 19444 24924 19445 24988
rect 19379 24923 19445 24924
rect 19382 20909 19442 24923
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 20483 22404 20549 22405
rect 20483 22340 20484 22404
rect 20548 22340 20549 22404
rect 20483 22339 20549 22340
rect 19379 20908 19445 20909
rect 19379 20844 19380 20908
rect 19444 20844 19445 20908
rect 19379 20843 19445 20844
rect 19563 19412 19629 19413
rect 19563 19348 19564 19412
rect 19628 19348 19629 19412
rect 19563 19347 19629 19348
rect 19566 10709 19626 19347
rect 19563 10708 19629 10709
rect 19563 10644 19564 10708
rect 19628 10644 19629 10708
rect 19563 10643 19629 10644
rect 18459 10164 18525 10165
rect 18459 10100 18460 10164
rect 18524 10100 18525 10164
rect 18459 10099 18525 10100
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17355 3636 17421 3637
rect 17355 3572 17356 3636
rect 17420 3572 17421 3636
rect 17355 3571 17421 3572
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 20486 1869 20546 22339
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 23427 19276 23493 19277
rect 23427 19212 23428 19276
rect 23492 19212 23493 19276
rect 23427 19211 23493 19212
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 21219 18052 21285 18053
rect 21219 17988 21220 18052
rect 21284 17988 21285 18052
rect 21219 17987 21285 17988
rect 21222 9621 21282 17987
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 21771 16692 21837 16693
rect 21771 16628 21772 16692
rect 21836 16628 21837 16692
rect 21771 16627 21837 16628
rect 21219 9620 21285 9621
rect 21219 9556 21220 9620
rect 21284 9556 21285 9620
rect 21219 9555 21285 9556
rect 21774 5541 21834 16627
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 21771 5540 21837 5541
rect 21771 5476 21772 5540
rect 21836 5476 21837 5540
rect 21771 5475 21837 5476
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 23430 4045 23490 19211
rect 23982 12069 24042 41379
rect 24715 18052 24781 18053
rect 24715 17988 24716 18052
rect 24780 17988 24781 18052
rect 24715 17987 24781 17988
rect 23979 12068 24045 12069
rect 23979 12004 23980 12068
rect 24044 12004 24045 12068
rect 23979 12003 24045 12004
rect 24718 4045 24778 17987
rect 23427 4044 23493 4045
rect 23427 3980 23428 4044
rect 23492 3980 23493 4044
rect 23427 3979 23493 3980
rect 24715 4044 24781 4045
rect 24715 3980 24716 4044
rect 24780 3980 24781 4044
rect 24715 3979 24781 3980
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 20483 1868 20549 1869
rect 20483 1804 20484 1868
rect 20548 1804 20549 1868
rect 20483 1803 20549 1804
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_
timestamp 1676037725
transform 1 0 11040 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1676037725
transform -1 0 18952 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _108_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1676037725
transform -1 0 22264 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _110_
timestamp 1676037725
transform -1 0 12604 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1676037725
transform -1 0 10580 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1676037725
transform -1 0 10672 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1676037725
transform -1 0 15732 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform -1 0 24932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 25024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1676037725
transform -1 0 22264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform -1 0 22264 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform -1 0 22264 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1676037725
transform -1 0 23000 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1676037725
transform -1 0 22264 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform -1 0 21068 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform -1 0 21896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1676037725
transform -1 0 22448 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform -1 0 21068 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform -1 0 21804 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform -1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform -1 0 20056 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform -1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform -1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1676037725
transform -1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform -1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform -1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform -1 0 18860 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform -1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform -1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform -1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform -1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform -1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 21804 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform -1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 23092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform -1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform -1 0 24932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform -1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform -1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1676037725
transform 1 0 5152 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 6532 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform -1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 9200 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 8280 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 9384 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 11408 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1676037725
transform 1 0 18400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1676037725
transform -1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform -1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform -1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1676037725
transform -1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform -1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1676037725
transform 1 0 14168 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform -1 0 21712 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform -1 0 25300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1676037725
transform -1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform -1 0 23092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform -1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1676037725
transform -1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1676037725
transform -1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform -1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1676037725
transform -1 0 24196 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1676037725
transform -1 0 25300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1676037725
transform -1 0 24288 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 11132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 14168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1676037725
transform -1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1676037725
transform -1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16928 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 15456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A0
timestamp 1676037725
transform -1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 14168 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1__S
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__S
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 15732 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__S
timestamp 1676037725
transform 1 0 14352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform -1 0 13892 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1__S
timestamp 1676037725
transform -1 0 12788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__S
timestamp 1676037725
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 17296 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__S
timestamp 1676037725
transform -1 0 15456 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform -1 0 11684 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 11040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 11684 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 10120 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 11316 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 8280 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 8832 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 15548 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform -1 0 16008 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 16928 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 19504 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform -1 0 25484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold5_A
timestamp 1676037725
transform -1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold10_A
timestamp 1676037725
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1676037725
transform -1 0 23184 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform -1 0 24564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform -1 0 24932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform -1 0 25576 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform -1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform -1 0 25576 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform -1 0 24840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform -1 0 25576 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform -1 0 24932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform -1 0 25576 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform -1 0 24932 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform -1 0 25576 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform -1 0 25576 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform -1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform -1 0 25576 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform -1 0 24840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform -1 0 25576 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform -1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform -1 0 25576 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform -1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform -1 0 25576 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform -1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform -1 0 25576 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform -1 0 24748 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform -1 0 24564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform -1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform -1 0 25576 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform -1 0 25576 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform -1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform -1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform -1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform -1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform -1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 5244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform -1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform -1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform -1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform -1 0 7636 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform -1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform -1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform -1 0 3680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform -1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform -1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform -1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform -1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform -1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform -1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform -1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform -1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform -1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform -1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform -1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform -1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform -1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform -1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform -1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform -1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform -1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform -1 0 13984 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform -1 0 15548 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform -1 0 17480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform -1 0 18308 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform -1 0 19136 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform -1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform -1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform -1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform -1 0 24196 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform -1 0 25576 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform -1 0 22816 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform -1 0 25208 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform -1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform -1 0 23552 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform -1 0 21436 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform -1 0 22724 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform -1 0 23368 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1676037725
transform -1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1676037725
transform -1 0 25208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1676037725
transform -1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1676037725
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1676037725
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22816 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23184 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22724 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24472 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23092 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 15456 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 11316 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15824 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15272 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15456 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24748 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 25576 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19688 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24472 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22356 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16744 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 16560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16744 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 7268 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__S
timestamp 1676037725
transform -1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 9016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform -1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18492 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15088 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 21620 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__A1
timestamp 1676037725
transform -1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1676037725
transform -1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 22448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l2_in_0__A0
timestamp 1676037725
transform -1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1676037725
transform -1 0 21712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_1__S
timestamp 1676037725
transform -1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8372 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 9108 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6440 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 9568 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8004 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform -1 0 10948 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform -1 0 9844 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 9384 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195
timestamp 1676037725
transform -1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform -1 0 8648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 9200 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13800 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform -1 0 12696 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13340 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13432 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform -1 0 13248 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform -1 0 11040 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196
timestamp 1676037725
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14720 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13800 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform -1 0 10856 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197
timestamp 1676037725
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17572 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform -1 0 16744 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 12512 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 10856 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9568 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 11224 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 13892 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 11592 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9384 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8924 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 10948 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 12696 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 10304 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform -1 0 8096 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform -1 0 8648 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 8464 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17756 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 11224 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 12604 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform -1 0 11224 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 12420 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform -1 0 18308 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform -1 0 15088 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform -1 0 15364 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform -1 0 15640 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform -1 0 16376 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform -1 0 21344 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 22172 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 19872 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 22080 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_247
timestamp 1676037725
transform 1 0 23828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_253
timestamp 1676037725
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1676037725
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_24
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1676037725
transform 1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_91
timestamp 1676037725
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1676037725
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1676037725
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1676037725
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_26
timestamp 1676037725
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1676037725
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1676037725
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_47 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_53
timestamp 1676037725
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1676037725
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_73
timestamp 1676037725
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_85
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1676037725
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1676037725
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_229
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_252
timestamp 1676037725
transform 1 0 24288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1676037725
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1676037725
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1676037725
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1676037725
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1676037725
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1676037725
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1676037725
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1676037725
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1676037725
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1676037725
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1676037725
transform 1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1676037725
transform 1 0 10580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1676037725
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_151
timestamp 1676037725
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1676037725
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1676037725
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1676037725
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_263
timestamp 1676037725
transform 1 0 25300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1676037725
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1676037725
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1676037725
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1676037725
transform 1 0 14536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1676037725
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_243
timestamp 1676037725
transform 1 0 23460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1676037725
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_130
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_180
timestamp 1676037725
transform 1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_253
timestamp 1676037725
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_258
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_129
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1676037725
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_150
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1676037725
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1676037725
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1676037725
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_130
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1676037725
transform 1 0 13616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1676037725
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_173
timestamp 1676037725
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1676037725
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_156
timestamp 1676037725
transform 1 0 15456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_169
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1676037725
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_248
timestamp 1676037725
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_118
timestamp 1676037725
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_126
timestamp 1676037725
transform 1 0 12696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_146
timestamp 1676037725
transform 1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1676037725
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_180
timestamp 1676037725
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_111
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_158
timestamp 1676037725
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_187
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1676037725
transform 1 0 22080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_262
timestamp 1676037725
transform 1 0 25208 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1676037725
transform 1 0 17112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1676037725
transform 1 0 19504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1676037725
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_265
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1676037725
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1676037725
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_155
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1676037725
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_174
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1676037725
transform 1 0 17848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1676037725
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_231
timestamp 1676037725
transform 1 0 22356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_235
timestamp 1676037725
transform 1 0 22724 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_131
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1676037725
transform 1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1676037725
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_236
timestamp 1676037725
transform 1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_263
timestamp 1676037725
transform 1 0 25300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1676037725
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1676037725
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1676037725
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_176
timestamp 1676037725
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1676037725
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_104
timestamp 1676037725
transform 1 0 10672 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1676037725
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_152
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_71
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1676037725
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_87
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1676037725
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1676037725
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1676037725
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1676037725
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1676037725
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_236
timestamp 1676037725
transform 1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1676037725
transform 1 0 24932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_263
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1676037725
transform 1 0 8372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1676037725
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1676037725
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_218
timestamp 1676037725
transform 1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_258
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1676037725
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_118
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1676037725
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1676037725
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1676037725
transform 1 0 20792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_230
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_263
timestamp 1676037725
transform 1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1676037725
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1676037725
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1676037725
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_164
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1676037725
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1676037725
transform 1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_107
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1676037725
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1676037725
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1676037725
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1676037725
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_100
timestamp 1676037725
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_150
timestamp 1676037725
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1676037725
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1676037725
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_264
timestamp 1676037725
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1676037725
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1676037725
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1676037725
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1676037725
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1676037725
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1676037725
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_108
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1676037725
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_190
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1676037725
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1676037725
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1676037725
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1676037725
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1676037725
transform 1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_228
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1676037725
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_143
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_155
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1676037725
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1676037725
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1676037725
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1676037725
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1676037725
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1676037725
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_95
timestamp 1676037725
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_110
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1676037725
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_158
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp 1676037725
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_230
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_259
timestamp 1676037725
transform 1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1676037725
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_118
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_148
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_154
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1676037725
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1676037725
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1676037725
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_248
timestamp 1676037725
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_259
timestamp 1676037725
transform 1 0 24932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1676037725
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1676037725
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_234
timestamp 1676037725
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_242
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_88
timestamp 1676037725
transform 1 0 9200 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1676037725
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1676037725
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1676037725
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1676037725
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_217
timestamp 1676037725
transform 1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1676037725
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1676037725
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1676037725
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_198
timestamp 1676037725
transform 1 0 19320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1676037725
transform 1 0 10212 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_117
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_127
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1676037725
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_183
timestamp 1676037725
transform 1 0 17940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1676037725
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1676037725
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1676037725
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1676037725
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_75
timestamp 1676037725
transform 1 0 8004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1676037725
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_100
timestamp 1676037725
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1676037725
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1676037725
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_195
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_201
timestamp 1676037725
transform 1 0 19596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_211
timestamp 1676037725
transform 1 0 20516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1676037725
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_96
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_100
timestamp 1676037725
transform 1 0 10304 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_108
timestamp 1676037725
transform 1 0 11040 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_119
timestamp 1676037725
transform 1 0 12052 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_143
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_146
timestamp 1676037725
transform 1 0 14536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_157
timestamp 1676037725
transform 1 0 15548 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_161
timestamp 1676037725
transform 1 0 15916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_181
timestamp 1676037725
transform 1 0 17756 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_216
timestamp 1676037725
transform 1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1676037725
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1676037725
transform 1 0 10212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1676037725
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1676037725
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_195
timestamp 1676037725
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_232
timestamp 1676037725
transform 1 0 22448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_238
timestamp 1676037725
transform 1 0 23000 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_107
timestamp 1676037725
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1676037725
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_143
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_155
timestamp 1676037725
transform 1 0 15364 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_219
timestamp 1676037725
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_258
timestamp 1676037725
transform 1 0 24840 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1676037725
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1676037725
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1676037725
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_199
timestamp 1676037725
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_242
timestamp 1676037725
transform 1 0 23368 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1676037725
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp 1676037725
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1676037725
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_152
timestamp 1676037725
transform 1 0 15088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_156
timestamp 1676037725
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1676037725
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_188
timestamp 1676037725
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_199
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1676037725
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1676037725
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_259
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_129
timestamp 1676037725
transform 1 0 12972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1676037725
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_174
timestamp 1676037725
transform 1 0 17112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_178
timestamp 1676037725
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_190
timestamp 1676037725
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_194
timestamp 1676037725
transform 1 0 18952 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_197
timestamp 1676037725
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1676037725
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_240
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1676037725
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_107
timestamp 1676037725
transform 1 0 10948 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_113
timestamp 1676037725
transform 1 0 11500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_125
timestamp 1676037725
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_152
timestamp 1676037725
transform 1 0 15088 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_156
timestamp 1676037725
transform 1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_167
timestamp 1676037725
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_185
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_219
timestamp 1676037725
transform 1 0 21252 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_223
timestamp 1676037725
transform 1 0 21620 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_229
timestamp 1676037725
transform 1 0 22172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_232
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1676037725
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_115
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_127
timestamp 1676037725
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1676037725
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1676037725
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp 1676037725
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_207
timestamp 1676037725
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1676037725
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_229
timestamp 1676037725
transform 1 0 22172 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1676037725
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_101
timestamp 1676037725
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_122
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_126
timestamp 1676037725
transform 1 0 12696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_162
timestamp 1676037725
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_168
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 1676037725
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_203
timestamp 1676037725
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1676037725
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_248
timestamp 1676037725
transform 1 0 23920 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp 1676037725
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1676037725
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_135
timestamp 1676037725
transform 1 0 13524 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_139
timestamp 1676037725
transform 1 0 13892 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1676037725
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_162
timestamp 1676037725
transform 1 0 16008 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_187
timestamp 1676037725
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_196
timestamp 1676037725
transform 1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_200
timestamp 1676037725
transform 1 0 19504 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_260
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1676037725
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1676037725
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_132
timestamp 1676037725
transform 1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_158
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp 1676037725
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1676037725
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1676037725
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1676037725
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_129
timestamp 1676037725
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1676037725
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_186
timestamp 1676037725
transform 1 0 18216 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_201
timestamp 1676037725
transform 1 0 19596 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_207
timestamp 1676037725
transform 1 0 20148 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1676037725
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_227
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1676037725
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1676037725
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_260
timestamp 1676037725
transform 1 0 25024 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_129
timestamp 1676037725
transform 1 0 12972 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_135
timestamp 1676037725
transform 1 0 13524 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_162
timestamp 1676037725
transform 1 0 16008 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1676037725
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1676037725
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1676037725
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1676037725
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_216
timestamp 1676037725
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1676037725
transform 1 0 22080 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_238
timestamp 1676037725
transform 1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_243
timestamp 1676037725
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_257
timestamp 1676037725
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_88
timestamp 1676037725
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_100
timestamp 1676037725
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1676037725
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_140
timestamp 1676037725
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_152
timestamp 1676037725
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_173
timestamp 1676037725
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_185
timestamp 1676037725
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_195
timestamp 1676037725
transform 1 0 19044 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 1676037725
transform 1 0 19780 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_213
timestamp 1676037725
transform 1 0 20700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 1676037725
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1676037725
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_90
timestamp 1676037725
transform 1 0 9384 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_102
timestamp 1676037725
transform 1 0 10488 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_114
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_126
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_155
timestamp 1676037725
transform 1 0 15364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_161
timestamp 1676037725
transform 1 0 15916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_169
timestamp 1676037725
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_190
timestamp 1676037725
transform 1 0 18584 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_205
timestamp 1676037725
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_237
timestamp 1676037725
transform 1 0 22908 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_241
timestamp 1676037725
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1676037725
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_154
timestamp 1676037725
transform 1 0 15272 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_160
timestamp 1676037725
transform 1 0 15824 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_171
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1676037725
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_201
timestamp 1676037725
transform 1 0 19596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_204
timestamp 1676037725
transform 1 0 19872 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_215
timestamp 1676037725
transform 1 0 20884 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1676037725
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1676037725
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1676037725
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_190
timestamp 1676037725
transform 1 0 18584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_219
timestamp 1676037725
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_232
timestamp 1676037725
transform 1 0 22448 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_236
timestamp 1676037725
transform 1 0 22816 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_174
timestamp 1676037725
transform 1 0 17112 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_186
timestamp 1676037725
transform 1 0 18216 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_194
timestamp 1676037725
transform 1 0 18952 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_215
timestamp 1676037725
transform 1 0 20884 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_219
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_263
timestamp 1676037725
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_166
timestamp 1676037725
transform 1 0 16376 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_174
timestamp 1676037725
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1676037725
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1676037725
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_202
timestamp 1676037725
transform 1 0 19688 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_215
timestamp 1676037725
transform 1 0 20884 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_227
timestamp 1676037725
transform 1 0 21988 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1676037725
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_220
timestamp 1676037725
transform 1 0 21344 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 1676037725
transform 1 0 24656 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1676037725
transform 1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1676037725
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1676037725
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1676037725
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1676037725
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1676037725
transform 1 0 15640 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_162
timestamp 1676037725
transform 1 0 16008 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_174
timestamp 1676037725
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1676037725
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1676037725
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_243
timestamp 1676037725
transform 1 0 23460 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1676037725
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_259
timestamp 1676037725
transform 1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1676037725
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_259
timestamp 1676037725
transform 1 0 24932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1676037725
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_117
timestamp 1676037725
transform 1 0 11868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_129
timestamp 1676037725
transform 1 0 12972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1676037725
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1676037725
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1676037725
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_236
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_248
timestamp 1676037725
transform 1 0 23920 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1676037725
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1676037725
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_257
timestamp 1676037725
transform 1 0 24748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1676037725
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_261
timestamp 1676037725
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 1676037725
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 1676037725
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_255
timestamp 1676037725
transform 1 0 24564 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_258
timestamp 1676037725
transform 1 0 24840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_259
timestamp 1676037725
transform 1 0 24932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_261
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_259
timestamp 1676037725
transform 1 0 24932 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1676037725
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_107
timestamp 1676037725
transform 1 0 10948 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_119
timestamp 1676037725
transform 1 0 12052 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 1676037725
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_89
timestamp 1676037725
transform 1 0 9292 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_117
timestamp 1676037725
transform 1 0 11868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_129
timestamp 1676037725
transform 1 0 12972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_141
timestamp 1676037725
transform 1 0 14076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_153
timestamp 1676037725
transform 1 0 15180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_165
timestamp 1676037725
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_100
timestamp 1676037725
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_112
timestamp 1676037725
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_124
timestamp 1676037725
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1676037725
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1676037725
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_257
timestamp 1676037725
transform 1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_229
timestamp 1676037725
transform 1 0 22172 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_261
timestamp 1676037725
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_101
timestamp 1676037725
transform 1 0 10396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1676037725
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_115
timestamp 1676037725
transform 1 0 11684 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_127
timestamp 1676037725
transform 1 0 12788 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_139
timestamp 1676037725
transform 1 0 13892 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_151
timestamp 1676037725
transform 1 0 14996 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_163
timestamp 1676037725
transform 1 0 16100 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_255
timestamp 1676037725
transform 1 0 24564 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_258
timestamp 1676037725
transform 1 0 24840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_107
timestamp 1676037725
transform 1 0 10948 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_113
timestamp 1676037725
transform 1 0 11500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_125
timestamp 1676037725
transform 1 0 12604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_137
timestamp 1676037725
transform 1 0 13708 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_157
timestamp 1676037725
transform 1 0 15548 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_179
timestamp 1676037725
transform 1 0 17572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_191
timestamp 1676037725
transform 1 0 18676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_147
timestamp 1676037725
transform 1 0 14628 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_159
timestamp 1676037725
transform 1 0 15732 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1676037725
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1676037725
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_129
timestamp 1676037725
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1676037725
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_170
timestamp 1676037725
transform 1 0 16744 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_182
timestamp 1676037725
transform 1 0 17848 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1676037725
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_259
timestamp 1676037725
transform 1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_99
timestamp 1676037725
transform 1 0 10212 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_106
timestamp 1676037725
transform 1 0 10856 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1676037725
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_121
timestamp 1676037725
transform 1 0 12236 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_127
timestamp 1676037725
transform 1 0 12788 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_160
timestamp 1676037725
transform 1 0 15824 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1676037725
transform 1 0 11500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_117
timestamp 1676037725
transform 1 0 11868 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1676037725
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1676037725
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1676037725
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_89
timestamp 1676037725
transform 1 0 9292 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_96
timestamp 1676037725
transform 1 0 9936 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_100
timestamp 1676037725
transform 1 0 10304 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_259
timestamp 1676037725
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1676037725
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_103
timestamp 1676037725
transform 1 0 10580 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_115
timestamp 1676037725
transform 1 0 11684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_127
timestamp 1676037725
transform 1 0 12788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_241
timestamp 1676037725
transform 1 0 23276 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_250
timestamp 1676037725
transform 1 0 24104 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_80
timestamp 1676037725
transform 1 0 8464 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_86
timestamp 1676037725
transform 1 0 9016 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_98
timestamp 1676037725
transform 1 0 10120 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_110
timestamp 1676037725
transform 1 0 11224 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_105
timestamp 1676037725
transform 1 0 10764 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_111
timestamp 1676037725
transform 1 0 11316 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_116
timestamp 1676037725
transform 1 0 11776 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_128
timestamp 1676037725
transform 1 0 12880 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1676037725
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1676037725
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_69
timestamp 1676037725
transform 1 0 7452 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_76
timestamp 1676037725
transform 1 0 8096 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_80
timestamp 1676037725
transform 1 0 8464 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_89
timestamp 1676037725
transform 1 0 9292 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_94
timestamp 1676037725
transform 1 0 9752 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_106
timestamp 1676037725
transform 1 0 10856 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1676037725
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_130
timestamp 1676037725
transform 1 0 13064 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_138
timestamp 1676037725
transform 1 0 13800 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1676037725
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1676037725
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1676037725
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_253
timestamp 1676037725
transform 1 0 24380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_256
timestamp 1676037725
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_69
timestamp 1676037725
transform 1 0 7452 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_74
timestamp 1676037725
transform 1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1676037725
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1676037725
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_103
timestamp 1676037725
transform 1 0 10580 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_115
timestamp 1676037725
transform 1 0 11684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1676037725
transform 1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_251
timestamp 1676037725
transform 1 0 24196 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_256
timestamp 1676037725
transform 1 0 24656 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1676037725
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_74
timestamp 1676037725
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_250
timestamp 1676037725
transform 1 0 24104 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_255
timestamp 1676037725
transform 1 0 24564 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1676037725
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1676037725
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1676037725
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_39
timestamp 1676037725
transform 1 0 4692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_43
timestamp 1676037725
transform 1 0 5060 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1676037725
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1676037725
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_233
timestamp 1676037725
transform 1 0 22540 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_236
timestamp 1676037725
transform 1 0 22816 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_244
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_250
timestamp 1676037725
transform 1 0 24104 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1676037725
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1676037725
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_47
timestamp 1676037725
transform 1 0 5428 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_59
timestamp 1676037725
transform 1 0 6532 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_76
timestamp 1676037725
transform 1 0 8096 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_229
timestamp 1676037725
transform 1 0 22172 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_234
timestamp 1676037725
transform 1 0 22632 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1676037725
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1676037725
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_89
timestamp 1676037725
transform 1 0 9292 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_106
timestamp 1676037725
transform 1 0 10856 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_136
timestamp 1676037725
transform 1 0 13616 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_146
timestamp 1676037725
transform 1 0 14536 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_153
timestamp 1676037725
transform 1 0 15180 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_157
timestamp 1676037725
transform 1 0 15548 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_174
timestamp 1676037725
transform 1 0 17112 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_178
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_187
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_209
timestamp 1676037725
transform 1 0 20332 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_221
timestamp 1676037725
transform 1 0 21436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_231
timestamp 1676037725
transform 1 0 22356 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_235
timestamp 1676037725
transform 1 0 22724 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_240
timestamp 1676037725
transform 1 0 23184 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1676037725
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25300 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform -1 0 24288 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform 1 0 24656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform -1 0 25300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1676037725
transform -1 0 24104 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1676037725
transform -1 0 24104 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1676037725
transform -1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1676037725
transform -1 0 25392 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1676037725
transform 1 0 24656 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 24380 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform -1 0 25392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform -1 0 25392 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform -1 0 25392 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform -1 0 25392 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform -1 0 25392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform -1 0 25392 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1676037725
transform -1 0 25392 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform -1 0 25392 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform -1 0 25392 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform -1 0 24104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform -1 0 24104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform -1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform -1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform -1 0 8648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform -1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform -1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform -1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform -1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform -1 0 11960 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform -1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform -1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform -1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1676037725
transform -1 0 6072 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 14260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform -1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25392 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform -1 0 25392 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1676037725
transform -1 0 25392 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25392 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform -1 0 22632 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform -1 0 24104 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform -1 0 24840 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform -1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform -1 0 21068 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform -1 0 22356 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform -1 0 24104 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18952 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform -1 0 3036 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform -1 0 16376 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform -1 0 24104 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform -1 0 23552 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform -1 0 24104 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform -1 0 25392 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform -1 0 24104 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform -1 0 24104 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform -1 0 11224 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform -1 0 24104 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform -1 0 24104 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform -1 0 22264 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform -1 0 23552 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform -1 0 13800 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform -1 0 20148 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform -1 0 18860 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform -1 0 13800 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform -1 0 20884 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform -1 0 23460 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 21712 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform -1 0 22724 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform -1 0 16744 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform -1 0 21528 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform -1 0 18400 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform -1 0 21712 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform -1 0 21528 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform -1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform -1 0 14444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform -1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform -1 0 17572 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform -1 0 18308 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform -1 0 18308 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform -1 0 3496 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform -1 0 5428 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform -1 0 6072 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform -1 0 8096 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform -1 0 8648 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 9384 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 10764 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 12144 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 25116 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23368 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21252 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 25024 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23920 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21712 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 19780 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 18860 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18584 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17388 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20700 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24104 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23460 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21344 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 20884 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20608 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 22172 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 15272 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 12328 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9292 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 13616 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 14904 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 14812 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 12696 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 11224 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 9936 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12328 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 14904 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12696 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 14352 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 13616 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 12236 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 10948 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 16376 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 17020 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18676 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 18216 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 15548 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21436 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24104 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23092 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 24472 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 23828 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 21344 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 20608 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform -1 0 20332 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 19136 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform -1 0 20332 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform -1 0 25392 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153
timestamp 1676037725
transform -1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160
timestamp 1676037725
transform -1 0 21528 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22172 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform -1 0 20056 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22632 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163
timestamp 1676037725
transform -1 0 22264 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199
timestamp 1676037725
transform -1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201
timestamp 1676037725
transform -1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202
timestamp 1676037725
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 18216 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17020 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154
timestamp 1676037725
transform -1 0 19964 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22356 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1676037725
transform -1 0 25392 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156
timestamp 1676037725
transform -1 0 25024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157
timestamp 1676037725
transform -1 0 21528 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158
timestamp 1676037725
transform -1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18768 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 15916 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161
timestamp 1676037725
transform -1 0 21528 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__164
timestamp 1676037725
transform -1 0 7452 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 8464 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform -1 0 12512 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17204 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15180 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform -1 0 10028 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform -1 0 12972 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17112 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform -1 0 16008 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform -1 0 16284 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform -1 0 11500 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform -1 0 14352 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17848 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15272 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform -1 0 12144 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__192
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform -1 0 15272 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15640 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__193
timestamp 1676037725
transform -1 0 9384 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform -1 0 9844 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform -1 0 12788 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17112 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform -1 0 7452 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform -1 0 10764 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 15272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform -1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform -1 0 12328 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1676037725
transform -1 0 13064 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15640 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18952 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1676037725
transform -1 0 13616 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15824 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15364 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__169
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18952 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform -1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18308 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform -1 0 11224 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__172
timestamp 1676037725
transform -1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform -1 0 13064 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform -1 0 12512 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15088 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 18492 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform -1 0 14628 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform -1 0 17296 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__175
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform -1 0 14536 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__176
timestamp 1676037725
transform -1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform -1 0 16560 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform -1 0 18308 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 21528 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform -1 0 18676 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__177
timestamp 1676037725
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform -1 0 16376 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17664 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__178
timestamp 1676037725
transform -1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform -1 0 13800 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 21804 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform -1 0 14168 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__179
timestamp 1676037725
transform -1 0 14720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 13800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform -1 0 15548 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__182
timestamp 1676037725
transform -1 0 16376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1676037725
transform -1 0 18952 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__184
timestamp 1676037725
transform -1 0 16928 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform -1 0 18860 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform -1 0 20424 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20516 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1676037725
transform -1 0 19596 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__185
timestamp 1676037725
transform -1 0 18952 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform -1 0 21528 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21252 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1676037725
transform -1 0 20424 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform -1 0 22264 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform -1 0 21528 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__187
timestamp 1676037725
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20332 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__188
timestamp 1676037725
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__189
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__190
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__191
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1676037725
transform -1 0 11868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 9890 29070 9890 29070 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9798 30906 9798 30906 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9338 42670 9338 42670 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 9062 34170 9062 34170 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8648 37978 8648 37978 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 9016 19278 9016 19278 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 13202 13872 13202 13872 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal2 9154 12988 9154 12988 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 6578 14484 6578 14484 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 7912 17714 7912 17714 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 9522 14926 9522 14926 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 10120 11662 10120 11662 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 8556 13362 8556 13362 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 8372 20366 8372 20366 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 10718 13838 10718 13838 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 11592 18190 11592 18190 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal2 7774 19822 7774 19822 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 10120 17714 10120 17714 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 10810 18666 10810 18666 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal2 10994 26044 10994 26044 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 13570 9146 13570 9146 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9108 19346 9108 19346 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8970 30702 8970 30702 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13846 9418 13846 9418 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14168 10234 14168 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13386 12206 13386 12206 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9614 12886 9614 12886 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11132 14994 11132 14994 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10994 12410 10994 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9660 12954 9660 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9936 12682 9936 12682 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9614 19346 9614 19346 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15042 8058 15042 8058 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7958 17578 7958 17578 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8786 30226 8786 30226 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13478 8874 13478 8874 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14996 9418 14996 9418 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13018 11152 13018 11152 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14352 14246 14352 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12742 9078 12742 9078 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12650 11016 12650 11016 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9798 11866 9798 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11500 13158 11500 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10028 17510 10028 17510 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal3 15594 12580 15594 12580 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9982 23018 9982 23018 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9292 33966 9292 33966 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15456 12886 15456 12886 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 14314 13478 14314 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 11866 12742 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11224 16626 11224 16626 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 13386 15555 13386 15555 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13018 14586 13018 14586 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10672 20366 10672 20366 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11086 20570 11086 20570 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11408 18870 11408 18870 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13570 15674 13570 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10442 26486 10442 26486 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 29274 9200 29274 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 14030 12580 14030 12580 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 13110 11611 13110 11611 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12328 15402 12328 15402 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10350 18496 10350 18496 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11546 21590 11546 21590 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11684 18428 11684 18428 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10856 18938 10856 18938 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 13570 23647 13570 23647 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 21658 10350 21658 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 10948 42262 10948 42262 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 10534 44166 10534 44166 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 10948 44268 10948 44268 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 16238 44778 16238 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 10626 43554 10626 43554 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal2 10350 48994 10350 48994 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 10396 49130 10396 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal2 16514 46104 16514 46104 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9200 47430 9200 47430 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 9200 44370 9200 44370 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 9568 50286 9568 50286 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 13938 46614 13938 46614 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 7590 51748 7590 51748 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 7912 46138 7912 46138 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 12788 45526 12788 45526 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25346 54128 25346 54128 0 ccff_head
rlabel metal2 1518 2064 1518 2064 0 ccff_head_0
rlabel metal3 25860 748 25860 748 0 ccff_tail
rlabel metal1 1426 53618 1426 53618 0 ccff_tail_0
rlabel metal1 24702 25466 24702 25466 0 chanx_right_in[0]
rlabel metal2 25346 34391 25346 34391 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal1 25116 36142 25116 36142 0 chanx_right_in[12]
rlabel metal2 25254 36703 25254 36703 0 chanx_right_in[13]
rlabel metal2 25254 37655 25254 37655 0 chanx_right_in[14]
rlabel via2 25346 38301 25346 38301 0 chanx_right_in[15]
rlabel metal2 25346 39253 25346 39253 0 chanx_right_in[16]
rlabel metal2 25530 40137 25530 40137 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25254 41565 25254 41565 0 chanx_right_in[19]
rlabel metal2 25346 26061 25346 26061 0 chanx_right_in[1]
rlabel metal2 25254 42483 25254 42483 0 chanx_right_in[20]
rlabel metal2 25254 43231 25254 43231 0 chanx_right_in[21]
rlabel metal2 25254 44183 25254 44183 0 chanx_right_in[22]
rlabel via2 25346 44829 25346 44829 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47447 25346 47447 0 chanx_right_in[26]
rlabel via2 25254 48093 25254 48093 0 chanx_right_in[27]
rlabel metal2 25254 49011 25254 49011 0 chanx_right_in[28]
rlabel via2 25346 49725 25346 49725 0 chanx_right_in[29]
rlabel metal2 23874 27013 23874 27013 0 chanx_right_in[2]
rlabel metal2 24518 28985 24518 28985 0 chanx_right_in[3]
rlabel metal1 23414 29580 23414 29580 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel via2 25530 30923 25530 30923 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal1 24840 33286 24840 33286 0 chanx_right_in[8]
rlabel metal2 25346 33677 25346 33677 0 chanx_right_in[9]
rlabel metal2 22218 2057 22218 2057 0 chanx_right_out[0]
rlabel metal2 25162 9129 25162 9129 0 chanx_right_out[10]
rlabel metal2 23322 10863 23322 10863 0 chanx_right_out[11]
rlabel metal1 23046 11628 23046 11628 0 chanx_right_out[12]
rlabel metal1 24150 12274 24150 12274 0 chanx_right_out[13]
rlabel metal3 25584 12988 25584 12988 0 chanx_right_out[14]
rlabel metal2 23414 13583 23414 13583 0 chanx_right_out[15]
rlabel metal1 24150 14450 24150 14450 0 chanx_right_out[16]
rlabel metal2 23322 15249 23322 15249 0 chanx_right_out[17]
rlabel metal2 24702 15589 24702 15589 0 chanx_right_out[18]
rlabel metal2 23874 16813 23874 16813 0 chanx_right_out[19]
rlabel metal2 22126 2125 22126 2125 0 chanx_right_out[1]
rlabel metal1 23322 17782 23322 17782 0 chanx_right_out[20]
rlabel metal1 24104 18326 24104 18326 0 chanx_right_out[21]
rlabel metal2 23874 19159 23874 19159 0 chanx_right_out[22]
rlabel metal2 24610 19261 24610 19261 0 chanx_right_out[23]
rlabel metal1 24380 20910 24380 20910 0 chanx_right_out[24]
rlabel metal3 24618 21964 24618 21964 0 chanx_right_out[25]
rlabel metal1 24150 23154 24150 23154 0 chanx_right_out[26]
rlabel metal2 24794 23069 24794 23069 0 chanx_right_out[27]
rlabel metal3 25124 24412 25124 24412 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal2 19090 6018 19090 6018 0 chanx_right_out[2]
rlabel metal2 22586 8687 22586 8687 0 chanx_right_out[3]
rlabel metal1 20654 6256 20654 6256 0 chanx_right_out[4]
rlabel metal2 23322 6239 23322 6239 0 chanx_right_out[5]
rlabel metal3 25630 6460 25630 6460 0 chanx_right_out[6]
rlabel metal1 23966 7310 23966 7310 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[9]
rlabel metal1 1794 2414 1794 2414 0 chany_bottom_in_0[0]
rlabel metal2 5520 1700 5520 1700 0 chany_bottom_in_0[10]
rlabel metal1 5658 3978 5658 3978 0 chany_bottom_in_0[11]
rlabel metal1 6210 3366 6210 3366 0 chany_bottom_in_0[12]
rlabel metal2 6670 1761 6670 1761 0 chany_bottom_in_0[13]
rlabel metal1 7084 3502 7084 3502 0 chany_bottom_in_0[14]
rlabel metal2 7406 1761 7406 1761 0 chany_bottom_in_0[15]
rlabel metal1 7820 3026 7820 3026 0 chany_bottom_in_0[16]
rlabel metal1 8418 2380 8418 2380 0 chany_bottom_in_0[17]
rlabel metal1 8694 3502 8694 3502 0 chany_bottom_in_0[18]
rlabel metal1 7130 2448 7130 2448 0 chany_bottom_in_0[19]
rlabel metal2 2254 2098 2254 2098 0 chany_bottom_in_0[1]
rlabel metal1 9154 4114 9154 4114 0 chany_bottom_in_0[20]
rlabel metal1 9476 3502 9476 3502 0 chany_bottom_in_0[21]
rlabel metal1 9568 2414 9568 2414 0 chany_bottom_in_0[22]
rlabel metal2 10350 1761 10350 1761 0 chany_bottom_in_0[23]
rlabel metal1 10442 3468 10442 3468 0 chany_bottom_in_0[24]
rlabel metal1 10350 2992 10350 2992 0 chany_bottom_in_0[25]
rlabel metal2 11454 1761 11454 1761 0 chany_bottom_in_0[26]
rlabel metal2 11822 1095 11822 1095 0 chany_bottom_in_0[27]
rlabel metal2 12006 748 12006 748 0 chany_bottom_in_0[28]
rlabel metal2 12558 2132 12558 2132 0 chany_bottom_in_0[29]
rlabel metal1 2392 3026 2392 3026 0 chany_bottom_in_0[2]
rlabel metal1 2484 2414 2484 2414 0 chany_bottom_in_0[3]
rlabel metal2 3358 1761 3358 1761 0 chany_bottom_in_0[4]
rlabel metal1 3496 3978 3496 3978 0 chany_bottom_in_0[5]
rlabel metal1 4002 3910 4002 3910 0 chany_bottom_in_0[6]
rlabel metal1 4416 3162 4416 3162 0 chany_bottom_in_0[7]
rlabel metal1 4462 3570 4462 3570 0 chany_bottom_in_0[8]
rlabel metal1 5750 3026 5750 3026 0 chany_bottom_in_0[9]
rlabel metal2 12926 1231 12926 1231 0 chany_bottom_out_0[0]
rlabel metal1 17756 3094 17756 3094 0 chany_bottom_out_0[10]
rlabel metal2 16974 1588 16974 1588 0 chany_bottom_out_0[11]
rlabel metal1 17480 4522 17480 4522 0 chany_bottom_out_0[12]
rlabel metal1 18814 3570 18814 3570 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal2 18446 1571 18446 1571 0 chany_bottom_out_0[15]
rlabel metal2 18814 2098 18814 2098 0 chany_bottom_out_0[16]
rlabel metal2 19182 1761 19182 1761 0 chany_bottom_out_0[17]
rlabel metal2 19550 1588 19550 1588 0 chany_bottom_out_0[18]
rlabel metal2 19918 1792 19918 1792 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal1 20792 3978 20792 3978 0 chany_bottom_out_0[20]
rlabel metal2 20654 1761 20654 1761 0 chany_bottom_out_0[21]
rlabel metal1 18768 3366 18768 3366 0 chany_bottom_out_0[22]
rlabel metal2 21390 1860 21390 1860 0 chany_bottom_out_0[23]
rlabel metal2 21758 1761 21758 1761 0 chany_bottom_out_0[24]
rlabel metal2 22126 1095 22126 1095 0 chany_bottom_out_0[25]
rlabel metal1 22540 8398 22540 8398 0 chany_bottom_out_0[26]
rlabel metal2 22862 1554 22862 1554 0 chany_bottom_out_0[27]
rlabel metal2 23230 1690 23230 1690 0 chany_bottom_out_0[28]
rlabel metal2 23598 1163 23598 1163 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14260 3434 14260 3434 0 chany_bottom_out_0[3]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal2 15134 1622 15134 1622 0 chany_bottom_out_0[6]
rlabel metal1 15502 3400 15502 3400 0 chany_bottom_out_0[7]
rlabel metal1 16468 2958 16468 2958 0 chany_bottom_out_0[8]
rlabel metal1 16652 4046 16652 4046 0 chany_bottom_out_0[9]
rlabel metal1 21758 32198 21758 32198 0 clknet_0_prog_clk
rlabel metal2 6854 14416 6854 14416 0 clknet_4_0_0_prog_clk
rlabel metal1 11454 42126 11454 42126 0 clknet_4_10_0_prog_clk
rlabel metal1 14398 31246 14398 31246 0 clknet_4_11_0_prog_clk
rlabel metal1 18906 20434 18906 20434 0 clknet_4_12_0_prog_clk
rlabel metal2 23322 21828 23322 21828 0 clknet_4_13_0_prog_clk
rlabel metal1 20792 32334 20792 32334 0 clknet_4_14_0_prog_clk
rlabel metal1 22770 43758 22770 43758 0 clknet_4_15_0_prog_clk
rlabel metal1 11868 13362 11868 13362 0 clknet_4_1_0_prog_clk
rlabel metal1 6624 18734 6624 18734 0 clknet_4_2_0_prog_clk
rlabel metal1 12604 20434 12604 20434 0 clknet_4_3_0_prog_clk
rlabel metal2 16882 13129 16882 13129 0 clknet_4_4_0_prog_clk
rlabel metal1 20286 7412 20286 7412 0 clknet_4_5_0_prog_clk
rlabel metal2 16974 21522 16974 21522 0 clknet_4_6_0_prog_clk
rlabel metal2 20286 18258 20286 18258 0 clknet_4_7_0_prog_clk
rlabel metal1 13386 29172 13386 29172 0 clknet_4_8_0_prog_clk
rlabel metal2 14858 27744 14858 27744 0 clknet_4_9_0_prog_clk
rlabel metal2 2438 55226 2438 55226 0 gfpga_pad_io_soc_dir[0]
rlabel metal1 4002 53618 4002 53618 0 gfpga_pad_io_soc_dir[1]
rlabel metal1 5152 54230 5152 54230 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6578 54920 6578 54920 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 13662 56236 13662 56236 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14996 54162 14996 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16836 54162 16836 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 17756 54162 17756 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal1 9614 54094 9614 54094 0 gfpga_pad_io_soc_out[1]
rlabel metal1 10718 53652 10718 53652 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12282 56236 12282 56236 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54162 19228 54162 0 isol_n
rlabel metal1 24242 48110 24242 48110 0 net1
rlabel metal1 23598 39270 23598 39270 0 net10
rlabel metal2 22126 22780 22126 22780 0 net100
rlabel metal1 23828 22202 23828 22202 0 net101
rlabel metal2 23966 23052 23966 23052 0 net102
rlabel metal1 22678 25228 22678 25228 0 net103
rlabel metal2 23966 25670 23966 25670 0 net104
rlabel metal2 15318 4896 15318 4896 0 net105
rlabel metal1 18975 3706 18975 3706 0 net106
rlabel metal1 13800 5882 13800 5882 0 net107
rlabel metal2 21988 8092 21988 8092 0 net108
rlabel metal2 22678 5882 22678 5882 0 net109
rlabel metal1 24242 40154 24242 40154 0 net11
rlabel metal1 24334 16082 24334 16082 0 net110
rlabel metal2 10258 5151 10258 5151 0 net111
rlabel metal2 14122 8330 14122 8330 0 net112
rlabel metal3 14536 12444 14536 12444 0 net113
rlabel metal2 19918 7582 19918 7582 0 net114
rlabel metal2 19458 6970 19458 6970 0 net115
rlabel metal1 19228 4590 19228 4590 0 net116
rlabel metal2 19550 6188 19550 6188 0 net117
rlabel metal2 18722 5542 18722 5542 0 net118
rlabel metal2 13754 5678 13754 5678 0 net119
rlabel metal1 25898 40902 25898 40902 0 net12
rlabel metal1 20746 3502 20746 3502 0 net120
rlabel metal2 20838 8364 20838 8364 0 net121
rlabel metal1 23414 2448 23414 2448 0 net122
rlabel metal3 21873 16660 21873 16660 0 net123
rlabel metal3 16560 20876 16560 20876 0 net124
rlabel metal1 21459 3094 21459 3094 0 net125
rlabel via1 22218 8789 22218 8789 0 net126
rlabel metal1 20654 5270 20654 5270 0 net127
rlabel metal1 23828 5202 23828 5202 0 net128
rlabel metal1 23782 2618 23782 2618 0 net129
rlabel metal3 24449 41412 24449 41412 0 net13
rlabel metal1 18354 5270 18354 5270 0 net130
rlabel metal2 22218 4199 22218 4199 0 net131
rlabel metal1 21758 7854 21758 7854 0 net132
rlabel metal1 23230 3162 23230 3162 0 net133
rlabel metal2 13478 3519 13478 3519 0 net134
rlabel metal1 14306 2618 14306 2618 0 net135
rlabel metal3 17319 15300 17319 15300 0 net136
rlabel metal1 14306 2414 14306 2414 0 net137
rlabel metal2 14858 5678 14858 5678 0 net138
rlabel metal1 16836 2414 16836 2414 0 net139
rlabel metal2 24702 24072 24702 24072 0 net14
rlabel metal2 17526 7004 17526 7004 0 net140
rlabel metal1 17434 13226 17434 13226 0 net141
rlabel metal1 18400 4114 18400 4114 0 net142
rlabel metal1 5106 53210 5106 53210 0 net143
rlabel metal1 5980 52666 5980 52666 0 net144
rlabel metal2 6026 52836 6026 52836 0 net145
rlabel metal2 9246 52564 9246 52564 0 net146
rlabel metal1 8372 51578 8372 51578 0 net147
rlabel metal2 9614 52326 9614 52326 0 net148
rlabel metal2 10718 51442 10718 51442 0 net149
rlabel metal1 23092 42534 23092 42534 0 net15
rlabel metal2 11730 51748 11730 51748 0 net150
rlabel metal1 18262 26010 18262 26010 0 net151
rlabel metal1 17940 27438 17940 27438 0 net152
rlabel metal2 24794 16524 24794 16524 0 net153
rlabel metal1 19872 28186 19872 28186 0 net154
rlabel metal1 22586 27098 22586 27098 0 net155
rlabel metal2 24978 28798 24978 28798 0 net156
rlabel metal1 21942 30226 21942 30226 0 net157
rlabel metal2 20286 30464 20286 30464 0 net158
rlabel metal2 19182 29376 19182 29376 0 net159
rlabel metal1 24702 43146 24702 43146 0 net16
rlabel metal1 22034 19346 22034 19346 0 net160
rlabel metal1 22080 17170 22080 17170 0 net161
rlabel metal1 19688 22746 19688 22746 0 net162
rlabel metal2 22218 21250 22218 21250 0 net163
rlabel metal1 7728 17306 7728 17306 0 net164
rlabel metal1 7222 12818 7222 12818 0 net165
rlabel metal2 8234 12546 8234 12546 0 net166
rlabel metal1 13478 17646 13478 17646 0 net167
rlabel metal2 13202 17408 13202 17408 0 net168
rlabel metal1 15364 16218 15364 16218 0 net169
rlabel metal1 25438 44166 25438 44166 0 net17
rlabel metal2 9982 21216 9982 21216 0 net170
rlabel metal2 12742 10914 12742 10914 0 net171
rlabel metal2 12650 7616 12650 7616 0 net172
rlabel metal1 15410 7854 15410 7854 0 net173
rlabel metal1 17296 14314 17296 14314 0 net174
rlabel metal1 14214 15130 14214 15130 0 net175
rlabel metal1 15916 16558 15916 16558 0 net176
rlabel metal2 15962 15232 15962 15232 0 net177
rlabel metal2 13386 8126 13386 8126 0 net178
rlabel metal1 15962 4454 15962 4454 0 net179
rlabel metal1 25116 40358 25116 40358 0 net18
rlabel metal1 18952 5678 18952 5678 0 net180
rlabel metal1 11408 21658 11408 21658 0 net181
rlabel metal2 21114 7582 21114 7582 0 net182
rlabel metal1 21574 9690 21574 9690 0 net183
rlabel metal2 18446 11968 18446 11968 0 net184
rlabel metal1 19044 12274 19044 12274 0 net185
rlabel metal2 20010 11390 20010 11390 0 net186
rlabel metal2 24610 6494 24610 6494 0 net187
rlabel metal2 11178 4403 11178 4403 0 net188
rlabel metal1 21114 2482 21114 2482 0 net189
rlabel metal2 25024 40732 25024 40732 0 net19
rlabel metal1 21252 3162 21252 3162 0 net190
rlabel metal1 11592 7854 11592 7854 0 net191
rlabel metal2 11730 19584 11730 19584 0 net192
rlabel metal2 9430 17408 9430 17408 0 net193
rlabel metal1 11270 12954 11270 12954 0 net194
rlabel metal2 11914 10302 11914 10302 0 net195
rlabel metal1 15410 23086 15410 23086 0 net196
rlabel metal1 16008 25874 16008 25874 0 net197
rlabel metal1 20332 21522 20332 21522 0 net198
rlabel metal1 24978 22032 24978 22032 0 net199
rlabel metal1 1794 4522 1794 4522 0 net2
rlabel metal1 24978 40902 24978 40902 0 net20
rlabel metal1 24380 24242 24380 24242 0 net200
rlabel metal1 20884 23154 20884 23154 0 net201
rlabel metal2 18538 24650 18538 24650 0 net202
rlabel metal1 24932 3366 24932 3366 0 net203
rlabel metal1 21574 43622 21574 43622 0 net204
rlabel metal2 25254 3706 25254 3706 0 net205
rlabel metal2 24610 2108 24610 2108 0 net206
rlabel metal1 24150 3706 24150 3706 0 net207
rlabel metal1 2622 3536 2622 3536 0 net208
rlabel metal1 5014 4522 5014 4522 0 net209
rlabel metal1 25944 33354 25944 33354 0 net21
rlabel metal2 24702 53754 24702 53754 0 net210
rlabel metal1 22632 47974 22632 47974 0 net211
rlabel metal1 2484 3910 2484 3910 0 net212
rlabel metal1 1794 3706 1794 3706 0 net213
rlabel metal1 24380 54162 24380 54162 0 net214
rlabel metal2 24610 52700 24610 52700 0 net215
rlabel metal1 25530 47974 25530 47974 0 net22
rlabel metal1 25392 49062 25392 49062 0 net23
rlabel metal2 25070 32164 25070 32164 0 net24
rlabel metal1 24886 20808 24886 20808 0 net25
rlabel metal1 24564 23086 24564 23086 0 net26
rlabel metal2 22494 27744 22494 27744 0 net27
rlabel metal1 23230 26350 23230 26350 0 net28
rlabel metal1 25116 26282 25116 26282 0 net29
rlabel metal2 19642 14144 19642 14144 0 net3
rlabel metal1 25116 31926 25116 31926 0 net30
rlabel metal1 25622 33286 25622 33286 0 net31
rlabel metal1 25714 33830 25714 33830 0 net32
rlabel metal2 7130 2040 7130 2040 0 net33
rlabel metal2 13846 14093 13846 14093 0 net34
rlabel metal1 12052 12614 12052 12614 0 net35
rlabel metal1 6624 3366 6624 3366 0 net36
rlabel metal2 6762 4658 6762 4658 0 net37
rlabel metal1 11270 12682 11270 12682 0 net38
rlabel metal1 12926 14926 12926 14926 0 net39
rlabel metal1 22770 34714 22770 34714 0 net4
rlabel metal2 14766 5916 14766 5916 0 net40
rlabel metal2 12190 12903 12190 12903 0 net41
rlabel metal2 8602 5746 8602 5746 0 net42
rlabel metal1 7912 2278 7912 2278 0 net43
rlabel metal1 7682 17170 7682 17170 0 net44
rlabel metal2 12466 6579 12466 6579 0 net45
rlabel metal1 14122 10574 14122 10574 0 net46
rlabel metal1 14766 9078 14766 9078 0 net47
rlabel metal2 17894 11594 17894 11594 0 net48
rlabel metal2 15318 10064 15318 10064 0 net49
rlabel metal1 25668 34918 25668 34918 0 net5
rlabel metal1 16514 9486 16514 9486 0 net50
rlabel metal1 18446 13430 18446 13430 0 net51
rlabel metal1 15732 9894 15732 9894 0 net52
rlabel metal1 16192 2346 16192 2346 0 net53
rlabel metal1 18354 10030 18354 10030 0 net54
rlabel metal1 2438 2924 2438 2924 0 net55
rlabel metal1 10534 21862 10534 21862 0 net56
rlabel metal1 11546 19686 11546 19686 0 net57
rlabel metal1 9062 17170 9062 17170 0 net58
rlabel metal1 7038 12716 7038 12716 0 net59
rlabel metal1 25990 36006 25990 36006 0 net6
rlabel metal1 8004 12818 8004 12818 0 net60
rlabel metal1 11822 17034 11822 17034 0 net61
rlabel metal1 13524 15334 13524 15334 0 net62
rlabel metal1 13524 53958 13524 53958 0 net63
rlabel metal2 13938 50286 13938 50286 0 net64
rlabel metal1 16790 46002 16790 46002 0 net65
rlabel metal1 17618 53958 17618 53958 0 net66
rlabel metal1 18262 54162 18262 54162 0 net67
rlabel metal2 7958 3417 7958 3417 0 net68
rlabel metal2 26312 35880 26312 35880 0 net69
rlabel metal1 25484 36550 25484 36550 0 net7
rlabel metal1 25852 51238 25852 51238 0 net70
rlabel metal1 16882 31960 16882 31960 0 net71
rlabel metal1 26036 51782 26036 51782 0 net72
rlabel metal1 22448 34374 22448 34374 0 net73
rlabel metal1 20378 32538 20378 32538 0 net74
rlabel metal1 24380 52870 24380 52870 0 net75
rlabel metal1 22494 32198 22494 32198 0 net76
rlabel metal2 16790 32980 16790 32980 0 net77
rlabel metal2 22264 35880 22264 35880 0 net78
rlabel metal1 23828 53414 23828 53414 0 net79
rlabel metal1 25576 37638 25576 37638 0 net8
rlabel metal1 19734 33014 19734 33014 0 net80
rlabel metal2 20424 14756 20424 14756 0 net81
rlabel metal2 5566 51986 5566 51986 0 net82
rlabel metal1 16330 6256 16330 6256 0 net83
rlabel metal1 15410 8500 15410 8500 0 net84
rlabel metal1 24334 7990 24334 7990 0 net85
rlabel metal1 24518 6426 24518 6426 0 net86
rlabel metal1 24564 11322 24564 11322 0 net87
rlabel metal1 25024 14246 25024 14246 0 net88
rlabel metal2 24058 13668 24058 13668 0 net89
rlabel metal1 25346 38182 25346 38182 0 net9
rlabel metal1 24564 13498 24564 13498 0 net90
rlabel metal1 22172 12954 22172 12954 0 net91
rlabel metal1 24380 12410 24380 12410 0 net92
rlabel metal1 22448 14042 22448 14042 0 net93
rlabel metal2 15778 3842 15778 3842 0 net94
rlabel metal1 24150 16762 24150 16762 0 net95
rlabel metal2 22218 18428 22218 18428 0 net96
rlabel metal2 22770 19482 22770 19482 0 net97
rlabel metal1 23736 18258 23736 18258 0 net98
rlabel metal1 21551 21046 21551 21046 0 net99
rlabel metal1 18354 24106 18354 24106 0 prog_clk
rlabel metal1 24518 4114 24518 4114 0 prog_reset
rlabel metal2 25254 50711 25254 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 25254 51323 25254 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 25254 52275 25254 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel via2 25530 52955 25530 52955 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 22586 53618 22586 53618 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 24932 53210 24932 53210 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25860 55420 25860 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 20562 56236 20562 56236 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21942 56236 21942 56236 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 23138 55711 23138 55711 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24288 52462 24288 52462 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 17066 44948 17066 44948 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21804 35258 21804 35258 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 21114 35615 21114 35615 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 24794 32742 24794 32742 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18722 14042 18722 14042 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal2 21666 19482 21666 19482 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal2 20194 18530 20194 18530 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 23092 21454 23092 21454 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal1 25392 24718 25392 24718 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 25024 23834 25024 23834 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 23000 27846 23000 27846 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 25162 27540 25162 27540 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 20240 26418 20240 26418 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal2 22126 28118 22126 28118 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal1 18354 26758 18354 26758 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal2 22586 27506 22586 27506 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal1 18354 30634 18354 30634 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal1 19550 29546 19550 29546 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal1 18170 31858 18170 31858 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 17112 31722 17112 31722 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 25162 19924 25162 19924 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal1 24288 20026 24288 20026 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 21068 31858 21068 31858 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal1 20240 31858 20240 31858 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal1 23644 30158 23644 30158 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 23322 31790 23322 31790 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 25346 32198 25346 32198 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal1 24886 32946 24886 32946 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 22908 34034 22908 34034 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal2 22310 34340 22310 34340 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 20010 33286 20010 33286 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel via1 22126 34170 22126 34170 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 19228 29070 19228 29070 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 21206 33150 21206 33150 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal2 23322 20298 23322 20298 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 25070 21454 25070 21454 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 23966 29070 23966 29070 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 19780 24038 19780 24038 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal1 21252 21862 21252 21862 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal2 22310 25568 22310 25568 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 11500 26554 11500 26554 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal1 18492 43622 18492 43622 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal1 8464 16762 8464 16762 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal1 11040 24038 11040 24038 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 8970 19142 8970 19142 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal1 14812 25330 14812 25330 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 6854 12784 6854 12784 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal1 10948 20026 10948 20026 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 8878 18938 8878 18938 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 14536 22066 14536 22066 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal1 12512 20774 12512 20774 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal2 14490 19822 14490 19822 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 12880 20366 12880 20366 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal2 11822 14824 11822 14824 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 12926 16626 12926 16626 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal2 11086 28322 11086 28322 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal2 13478 27744 13478 27744 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal1 12995 27506 12995 27506 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 12466 10540 12466 10540 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal1 10488 11186 10488 11186 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal2 10810 6460 10810 6460 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal2 9338 8058 9338 8058 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal1 12650 6834 12650 6834 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 11454 6222 11454 6222 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal1 16330 14450 16330 14450 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel metal2 14076 12750 14076 12750 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 16330 20026 16330 20026 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 14720 19754 14720 19754 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal1 18124 20366 18124 20366 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 15548 20774 15548 20774 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal1 18492 18054 18492 18054 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 17066 18190 17066 18190 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal1 16606 11254 16606 11254 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal2 16422 17238 16422 17238 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal1 16192 4998 16192 4998 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal2 13570 6698 13570 6698 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16737 5882 16737 5882 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15410 5134 15410 5134 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 13294 28390 13294 28390 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal1 13064 30158 13064 30158 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 13478 29036 13478 29036 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal2 21298 7038 21298 7038 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal1 17250 6698 17250 6698 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal2 21298 11424 21298 11424 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal1 19504 9146 19504 9146 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 20516 15334 20516 15334 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal1 19688 15402 19688 15402 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal1 20930 15980 20930 15980 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 21942 16592 21942 16592 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal1 21666 14416 21666 14416 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal1 22218 15538 22218 15538 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal2 24150 10030 24150 10030 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal1 20930 12716 20930 12716 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal1 23690 7990 23690 7990 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal1 22632 7922 22632 7922 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal1 20700 5134 20700 5134 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal1 21850 6426 21850 6426 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 18630 7514 18630 7514 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal1 19320 7310 19320 7310 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 17243 13702 17243 13702 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal2 13754 24548 13754 24548 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal2 15134 28152 15134 28152 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal1 11914 24106 11914 24106 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal2 16238 26962 16238 26962 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal2 9384 18428 9384 18428 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal1 15640 7718 15640 7718 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20654 19482 20654 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20470 20400 20470 20400 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 15062 19458 15062 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21344 15130 21344 15130 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 25162 21998 25162 21998 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 15028 21022 15028 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19596 16422 19596 16422 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 22632 24786 22632 24786 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21344 18156 21344 18156 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18906 15878 18906 15878 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal1 21436 23834 21436 23834 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19918 20876 19918 20876 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17250 15946 17250 15946 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 18860 24174 18860 24174 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18492 16150 18492 16150 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16744 17646 16744 17646 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 18630 25942 18630 25942 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 17714 17158 17714 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14352 6630 14352 6630 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 17802 27302 17802 27302 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 19346 16284 19346 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16238 7990 16238 7990 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal2 25070 19244 25070 19244 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22264 10642 22264 10642 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13800 12070 13800 12070 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal2 21666 30022 21666 30022 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19228 19822 19228 19822 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 21183 18020 21183 18020 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 22954 31926 22954 31926 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21298 22542 21298 22542 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19964 9962 19964 9962 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 25300 32742 25300 32742 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21482 18700 21482 18700 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 19665 19380 19665 19380 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal1 22632 30294 22632 30294 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21896 30022 21896 30022 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19044 16388 19044 16388 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal1 21298 35530 21298 35530 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19734 20502 19734 20502 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11040 12886 11040 12886 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 19872 35530 19872 35530 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17296 21590 17296 21590 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21114 13838 21114 13838 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 23368 19482 23368 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21114 13940 21114 13940 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16744 12614 16744 12614 0 sb_0__8_.mux_bottom_track_51.out
rlabel metal1 23460 17306 23460 17306 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 12852 20194 12852 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15916 15436 15916 15436 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal1 20010 22984 20010 22984 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20102 23086 20102 23086 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 17238 18308 17238 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17526 8840 17526 8840 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22540 21658 22540 21658 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel viali 20470 14380 20470 14380 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21574 25364 21574 25364 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 14122 32742 14122 32742 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14076 31926 14076 31926 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12006 26894 12006 26894 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10120 16966 10120 16966 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12972 24650 12972 24650 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15226 20230 15226 20230 0 sb_0__8_.mux_right_track_10.out
rlabel metal2 11730 24310 11730 24310 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11638 24786 11638 24786 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10764 18326 10764 18326 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8970 18054 8970 18054 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 15042 18734 15042 18734 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16882 20026 16882 20026 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 12236 18802 12236 18802 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11546 18666 11546 18666 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14582 19414 14582 19414 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21666 20944 21666 20944 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 15456 22134 15456 22134 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13524 17850 13524 17850 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15732 21862 15732 21862 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22034 18768 22034 18768 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 15364 20570 15364 20570 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14490 17306 14490 17306 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18998 19380 18998 19380 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21850 16456 21850 16456 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 14720 16218 14720 16218 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17664 16558 17664 16558 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 25296 20838 25296 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 13662 27438 13662 27438 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13662 27370 13662 27370 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12558 26010 12558 26010 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 9982 23766 9982 23766 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 16882 25942 16882 25942 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18262 12920 18262 12920 0 sb_0__8_.mux_right_track_20.out
rlabel metal2 12650 11016 12650 11016 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18216 12818 18216 12818 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 10778 21482 10778 0 sb_0__8_.mux_right_track_22.out
rlabel metal2 12558 6732 12558 6732 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14950 7514 14950 7514 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18722 10506 18722 10506 0 sb_0__8_.mux_right_track_24.out
rlabel metal1 12558 6086 12558 6086 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16422 7990 16422 7990 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21206 13736 21206 13736 0 sb_0__8_.mux_right_track_26.out
rlabel metal2 14582 13226 14582 13226 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20194 14076 20194 14076 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 17544 20838 17544 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 17020 23494 17020 23494 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14490 15096 14490 15096 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20654 17612 20654 17612 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23230 17374 23230 17374 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 18078 19822 18078 19822 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16514 18054 16514 18054 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21252 17646 21252 17646 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22310 15606 22310 15606 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 19596 17646 19596 17646 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16330 16354 16330 16354 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21666 15504 21666 15504 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21758 8534 21758 8534 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 17572 18598 17572 18598 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13754 7752 13754 7752 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21528 11118 21528 11118 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13662 6681 13662 6681 0 sb_0__8_.mux_right_track_36.out
rlabel metal1 15732 6426 15732 6426 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15778 6154 15778 6154 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15916 3978 15916 3978 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 17066 5746 17066 5746 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16790 4114 16790 4114 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 25160 17802 25160 0 sb_0__8_.mux_right_track_4.out
rlabel metal2 16054 29376 16054 29376 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15962 29648 15962 29648 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14260 25874 14260 25874 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 11454 23902 11454 23902 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 17618 25500 17618 25500 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 10626 4828 10626 4828 0 sb_0__8_.mux_right_track_40.out
rlabel metal1 20930 7514 20930 7514 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20930 6137 20930 6137 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18906 5117 18906 5117 0 sb_0__8_.mux_right_track_42.out
rlabel metal1 20930 10574 20930 10574 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19090 10574 19090 10574 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 16014 24564 16014 0 sb_0__8_.mux_right_track_44.out
rlabel metal2 19918 17952 19918 17952 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 14994 19458 14994 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21620 14858 21620 14858 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 12926 5219 12926 5219 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 20424 21862 20424 21862 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19780 12954 19780 12954 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 15776 21482 15776 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23276 13226 23276 13226 0 sb_0__8_.mux_right_track_48.out
rlabel metal2 21758 17340 21758 17340 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21160 14246 21160 14246 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23092 14246 23092 14246 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13570 5644 13570 5644 0 sb_0__8_.mux_right_track_50.out
rlabel metal2 21482 12517 21482 12517 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17342 6324 17342 6324 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 2618 18814 2618 0 sb_0__8_.mux_right_track_52.out
rlabel metal1 23644 9962 23644 9962 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18998 2414 18998 2414 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8832 2550 8832 2550 0 sb_0__8_.mux_right_track_54.out
rlabel metal2 21022 5406 21022 5406 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20562 2958 20562 2958 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12650 5270 12650 5270 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 18078 7514 18078 7514 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13386 4624 13386 4624 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24794 7242 24794 7242 0 sb_0__8_.mux_right_track_58.out
rlabel metal2 17158 15232 17158 15232 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 17043 12580 17043 12580 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17618 13226 17618 13226 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22034 21971 22034 21971 0 sb_0__8_.mux_right_track_6.out
rlabel metal2 15778 28016 15778 28016 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 27098 16284 27098 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 23834 14904 23834 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 20026 12742 20026 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18078 23630 18078 23630 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17066 22712 17066 22712 0 sb_0__8_.mux_right_track_8.out
rlabel metal1 13616 23630 13616 23630 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13662 25160 13662 25160 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 22814 12558 22814 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10442 17306 10442 17306 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13340 21862 13340 21862 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
