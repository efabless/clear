magic
tech sky130A
magscale 1 2
timestamp 1656240995
<< viali >>
rect 5733 14569 5767 14603
rect 6561 14569 6595 14603
rect 7665 14569 7699 14603
rect 10149 14569 10183 14603
rect 12357 14569 12391 14603
rect 14565 14569 14599 14603
rect 6929 14501 6963 14535
rect 14381 14501 14415 14535
rect 15117 14501 15151 14535
rect 15577 14501 15611 14535
rect 2237 14433 2271 14467
rect 3157 14433 3191 14467
rect 5181 14433 5215 14467
rect 6745 14433 6779 14467
rect 14933 14433 14967 14467
rect 1961 14365 1995 14399
rect 2881 14365 2915 14399
rect 4353 14365 4387 14399
rect 4629 14365 4663 14399
rect 4721 14365 4755 14399
rect 5917 14365 5951 14399
rect 7849 14365 7883 14399
rect 10333 14365 10367 14399
rect 12541 14365 12575 14399
rect 14749 14365 14783 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 16405 14365 16439 14399
rect 16773 14365 16807 14399
rect 17049 14365 17083 14399
rect 17693 14365 17727 14399
rect 17969 14365 18003 14399
rect 3433 14297 3467 14331
rect 6377 14297 6411 14331
rect 15301 14297 15335 14331
rect 16037 14297 16071 14331
rect 3341 14229 3375 14263
rect 4905 14229 4939 14263
rect 4997 14229 5031 14263
rect 5365 14229 5399 14263
rect 6009 14229 6043 14263
rect 8033 14229 8067 14263
rect 15945 14229 15979 14263
rect 16313 14229 16347 14263
rect 4169 14025 4203 14059
rect 4537 14025 4571 14059
rect 4997 14025 5031 14059
rect 5365 14025 5399 14059
rect 5457 14025 5491 14059
rect 6009 14025 6043 14059
rect 6929 14025 6963 14059
rect 12817 14025 12851 14059
rect 17417 14025 17451 14059
rect 7113 13957 7147 13991
rect 13231 13957 13265 13991
rect 15025 13957 15059 13991
rect 15761 13957 15795 13991
rect 17141 13957 17175 13991
rect 17509 13957 17543 13991
rect 2237 13889 2271 13923
rect 3341 13889 3375 13923
rect 3709 13889 3743 13923
rect 6377 13889 6411 13923
rect 10517 13889 10551 13923
rect 13001 13889 13035 13923
rect 13128 13889 13162 13923
rect 15209 13889 15243 13923
rect 15485 13889 15519 13923
rect 15945 13889 15979 13923
rect 16129 13889 16163 13923
rect 16405 13889 16439 13923
rect 16681 13889 16715 13923
rect 1961 13821 1995 13855
rect 2881 13821 2915 13855
rect 3157 13821 3191 13855
rect 3525 13821 3559 13855
rect 3893 13821 3927 13855
rect 4629 13821 4663 13855
rect 4721 13821 4755 13855
rect 5641 13821 5675 13855
rect 5825 13821 5859 13855
rect 10977 13821 11011 13855
rect 13553 13821 13587 13855
rect 16221 13821 16255 13855
rect 16957 13821 16991 13855
rect 17693 13821 17727 13855
rect 17969 13821 18003 13855
rect 3985 13753 4019 13787
rect 6561 13753 6595 13787
rect 15301 13753 15335 13787
rect 16865 13753 16899 13787
rect 6745 13685 6779 13719
rect 10793 13685 10827 13719
rect 3617 13481 3651 13515
rect 6837 13481 6871 13515
rect 1961 13345 1995 13379
rect 3065 13345 3099 13379
rect 5089 13345 5123 13379
rect 5917 13345 5951 13379
rect 7573 13345 7607 13379
rect 15025 13345 15059 13379
rect 17969 13345 18003 13379
rect 2237 13277 2271 13311
rect 3157 13277 3191 13311
rect 3801 13277 3835 13311
rect 5733 13277 5767 13311
rect 6469 13277 6503 13311
rect 7389 13277 7423 13311
rect 15117 13277 15151 13311
rect 17325 13277 17359 13311
rect 17693 13277 17727 13311
rect 2421 13209 2455 13243
rect 4169 13209 4203 13243
rect 4445 13209 4479 13243
rect 4905 13209 4939 13243
rect 5825 13209 5859 13243
rect 6653 13209 6687 13243
rect 15301 13209 15335 13243
rect 16957 13209 16991 13243
rect 17509 13209 17543 13243
rect 2513 13141 2547 13175
rect 2697 13141 2731 13175
rect 3249 13141 3283 13175
rect 3985 13141 4019 13175
rect 4537 13141 4571 13175
rect 4997 13141 5031 13175
rect 5365 13141 5399 13175
rect 6377 13141 6411 13175
rect 7021 13141 7055 13175
rect 7481 13141 7515 13175
rect 7941 13141 7975 13175
rect 17233 13141 17267 13175
rect 3525 12937 3559 12971
rect 3893 12937 3927 12971
rect 4537 12937 4571 12971
rect 4629 12937 4663 12971
rect 6193 12937 6227 12971
rect 6745 12937 6779 12971
rect 7297 12937 7331 12971
rect 7665 12937 7699 12971
rect 8585 12937 8619 12971
rect 15761 12937 15795 12971
rect 6653 12869 6687 12903
rect 8125 12869 8159 12903
rect 13461 12869 13495 12903
rect 16129 12869 16163 12903
rect 2697 12801 2731 12835
rect 3341 12801 3375 12835
rect 5365 12801 5399 12835
rect 5825 12801 5859 12835
rect 7757 12801 7791 12835
rect 8493 12801 8527 12835
rect 13369 12801 13403 12835
rect 13829 12801 13863 12835
rect 16313 12801 16347 12835
rect 16773 12801 16807 12835
rect 16957 12801 16991 12835
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 2421 12733 2455 12767
rect 2605 12733 2639 12767
rect 4721 12733 4755 12767
rect 5549 12733 5583 12767
rect 5733 12733 5767 12767
rect 6561 12733 6595 12767
rect 7849 12733 7883 12767
rect 9321 12733 9355 12767
rect 13645 12733 13679 12767
rect 15945 12733 15979 12767
rect 17693 12733 17727 12767
rect 17969 12733 18003 12767
rect 3157 12665 3191 12699
rect 9873 12665 9907 12699
rect 3065 12597 3099 12631
rect 3709 12597 3743 12631
rect 4169 12597 4203 12631
rect 4997 12597 5031 12631
rect 7113 12597 7147 12631
rect 9689 12597 9723 12631
rect 13001 12597 13035 12631
rect 16405 12597 16439 12631
rect 17141 12597 17175 12631
rect 17417 12597 17451 12631
rect 17601 12597 17635 12631
rect 2513 12393 2547 12427
rect 10701 12393 10735 12427
rect 13737 12393 13771 12427
rect 15025 12393 15059 12427
rect 8125 12325 8159 12359
rect 3525 12257 3559 12291
rect 4353 12257 4387 12291
rect 4721 12257 4755 12291
rect 4905 12257 4939 12291
rect 6009 12257 6043 12291
rect 6653 12257 6687 12291
rect 7849 12257 7883 12291
rect 9597 12257 9631 12291
rect 10333 12257 10367 12291
rect 12541 12257 12575 12291
rect 12909 12257 12943 12291
rect 14657 12257 14691 12291
rect 17325 12257 17359 12291
rect 17509 12257 17543 12291
rect 1961 12189 1995 12223
rect 2237 12189 2271 12223
rect 3249 12189 3283 12223
rect 4997 12189 5031 12223
rect 5825 12189 5859 12223
rect 6837 12189 6871 12223
rect 7757 12189 7791 12223
rect 9321 12189 9355 12223
rect 10241 12189 10275 12223
rect 13185 12189 13219 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 16313 12189 16347 12223
rect 17693 12189 17727 12223
rect 17969 12189 18003 12223
rect 2421 12121 2455 12155
rect 6745 12121 6779 12155
rect 10149 12121 10183 12155
rect 12449 12121 12483 12155
rect 13093 12121 13127 12155
rect 16497 12121 16531 12155
rect 2789 12053 2823 12087
rect 2881 12053 2915 12087
rect 3341 12053 3375 12087
rect 3801 12053 3835 12087
rect 4169 12053 4203 12087
rect 4261 12053 4295 12087
rect 5365 12053 5399 12087
rect 5457 12053 5491 12087
rect 5917 12053 5951 12087
rect 6285 12053 6319 12087
rect 7205 12053 7239 12087
rect 7297 12053 7331 12087
rect 7665 12053 7699 12087
rect 8953 12053 8987 12087
rect 9413 12053 9447 12087
rect 9781 12053 9815 12087
rect 11805 12053 11839 12087
rect 11989 12053 12023 12087
rect 12357 12053 12391 12087
rect 13553 12053 13587 12087
rect 13829 12053 13863 12087
rect 14105 12053 14139 12087
rect 15945 12053 15979 12087
rect 16037 12053 16071 12087
rect 16589 12053 16623 12087
rect 16865 12053 16899 12087
rect 17233 12053 17267 12087
rect 2605 11849 2639 11883
rect 2973 11849 3007 11883
rect 4077 11849 4111 11883
rect 4905 11849 4939 11883
rect 5457 11849 5491 11883
rect 5549 11849 5583 11883
rect 6469 11849 6503 11883
rect 7297 11849 7331 11883
rect 7757 11849 7791 11883
rect 8493 11849 8527 11883
rect 8585 11849 8619 11883
rect 10793 11849 10827 11883
rect 15761 11849 15795 11883
rect 17141 11849 17175 11883
rect 10149 11781 10183 11815
rect 10701 11781 10735 11815
rect 11897 11781 11931 11815
rect 15301 11781 15335 11815
rect 1501 11713 1535 11747
rect 2145 11713 2179 11747
rect 3433 11713 3467 11747
rect 3893 11713 3927 11747
rect 4445 11713 4479 11747
rect 6653 11713 6687 11747
rect 7665 11713 7699 11747
rect 9321 11713 9355 11747
rect 13461 11713 13495 11747
rect 13921 11713 13955 11747
rect 15209 11713 15243 11747
rect 15945 11713 15979 11747
rect 17049 11713 17083 11747
rect 17601 11713 17635 11747
rect 18061 11713 18095 11747
rect 18429 11713 18463 11747
rect 1961 11645 1995 11679
rect 2053 11645 2087 11679
rect 3065 11645 3099 11679
rect 3249 11645 3283 11679
rect 4537 11645 4571 11679
rect 4721 11645 4755 11679
rect 5365 11645 5399 11679
rect 7021 11645 7055 11679
rect 7849 11645 7883 11679
rect 8769 11645 8803 11679
rect 9413 11645 9447 11679
rect 9505 11645 9539 11679
rect 10977 11645 11011 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 15117 11645 15151 11679
rect 16405 11645 16439 11679
rect 17233 11645 17267 11679
rect 2513 11577 2547 11611
rect 3709 11577 3743 11611
rect 8953 11577 8987 11611
rect 14565 11577 14599 11611
rect 17785 11577 17819 11611
rect 1593 11509 1627 11543
rect 3617 11509 3651 11543
rect 5917 11509 5951 11543
rect 6193 11509 6227 11543
rect 6837 11509 6871 11543
rect 8125 11509 8159 11543
rect 9781 11509 9815 11543
rect 10333 11509 10367 11543
rect 11529 11509 11563 11543
rect 13093 11509 13127 11543
rect 14749 11509 14783 11543
rect 15669 11509 15703 11543
rect 16129 11509 16163 11543
rect 16313 11509 16347 11543
rect 16681 11509 16715 11543
rect 17969 11509 18003 11543
rect 18337 11509 18371 11543
rect 3525 11305 3559 11339
rect 4537 11305 4571 11339
rect 8769 11305 8803 11339
rect 15025 11305 15059 11339
rect 16865 11305 16899 11339
rect 2329 11237 2363 11271
rect 3433 11237 3467 11271
rect 5549 11237 5583 11271
rect 6377 11237 6411 11271
rect 9321 11237 9355 11271
rect 10977 11237 11011 11271
rect 14105 11237 14139 11271
rect 16589 11237 16623 11271
rect 2789 11169 2823 11203
rect 3893 11169 3927 11203
rect 4077 11169 4111 11203
rect 4813 11169 4847 11203
rect 6009 11169 6043 11203
rect 6193 11169 6227 11203
rect 6929 11169 6963 11203
rect 7757 11169 7791 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 9873 11169 9907 11203
rect 10793 11169 10827 11203
rect 11529 11169 11563 11203
rect 12909 11169 12943 11203
rect 13001 11169 13035 11203
rect 13553 11169 13587 11203
rect 14657 11169 14691 11203
rect 15761 11169 15795 11203
rect 17325 11169 17359 11203
rect 17509 11169 17543 11203
rect 1961 11101 1995 11135
rect 2237 11101 2271 11135
rect 2513 11101 2547 11135
rect 3065 11101 3099 11135
rect 4997 11101 5031 11135
rect 5917 11101 5951 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7573 11101 7607 11135
rect 8401 11101 8435 11135
rect 9689 11101 9723 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 13093 11101 13127 11135
rect 14565 11101 14599 11135
rect 15485 11101 15519 11135
rect 16221 11101 16255 11135
rect 16313 11101 16347 11135
rect 16773 11101 16807 11135
rect 17693 11101 17727 11135
rect 17969 11101 18003 11135
rect 2973 11033 3007 11067
rect 4905 11033 4939 11067
rect 7665 11033 7699 11067
rect 11345 11033 11379 11067
rect 13829 11033 13863 11067
rect 14473 11033 14507 11067
rect 15577 11033 15611 11067
rect 4169 10965 4203 10999
rect 5365 10965 5399 10999
rect 7205 10965 7239 10999
rect 8953 10965 8987 10999
rect 9229 10965 9263 10999
rect 9781 10965 9815 10999
rect 10149 10965 10183 10999
rect 11437 10965 11471 10999
rect 13461 10965 13495 10999
rect 15117 10965 15151 10999
rect 16037 10965 16071 10999
rect 16497 10965 16531 10999
rect 17233 10965 17267 10999
rect 2053 10761 2087 10795
rect 2513 10761 2547 10795
rect 2697 10761 2731 10795
rect 3065 10761 3099 10795
rect 3617 10761 3651 10795
rect 4077 10761 4111 10795
rect 4261 10761 4295 10795
rect 5825 10761 5859 10795
rect 5917 10761 5951 10795
rect 12909 10761 12943 10795
rect 13277 10761 13311 10795
rect 14473 10761 14507 10795
rect 15209 10761 15243 10795
rect 15761 10761 15795 10795
rect 16221 10761 16255 10795
rect 16681 10761 16715 10795
rect 17509 10761 17543 10795
rect 3709 10693 3743 10727
rect 3893 10693 3927 10727
rect 4629 10693 4663 10727
rect 6929 10693 6963 10727
rect 14381 10693 14415 10727
rect 1593 10625 1627 10659
rect 3157 10625 3191 10659
rect 5273 10625 5307 10659
rect 6561 10625 6595 10659
rect 6745 10625 6779 10659
rect 7389 10625 7423 10659
rect 8217 10625 8251 10659
rect 9597 10625 9631 10659
rect 10517 10625 10551 10659
rect 11345 10625 11379 10659
rect 11897 10625 11931 10659
rect 13369 10625 13403 10659
rect 15301 10625 15335 10659
rect 16129 10625 16163 10659
rect 17049 10625 17083 10659
rect 18061 10625 18095 10659
rect 18429 10625 18463 10659
rect 1777 10557 1811 10591
rect 1961 10557 1995 10591
rect 3341 10557 3375 10591
rect 4721 10557 4755 10591
rect 4813 10557 4847 10591
rect 6101 10557 6135 10591
rect 7481 10557 7515 10591
rect 7665 10557 7699 10591
rect 8309 10557 8343 10591
rect 8493 10557 8527 10591
rect 8677 10557 8711 10591
rect 8953 10557 8987 10591
rect 10609 10557 10643 10591
rect 10793 10557 10827 10591
rect 11713 10557 11747 10591
rect 11805 10557 11839 10591
rect 12449 10557 12483 10591
rect 13461 10557 13495 10591
rect 14565 10557 14599 10591
rect 15393 10557 15427 10591
rect 16313 10557 16347 10591
rect 17141 10557 17175 10591
rect 17325 10557 17359 10591
rect 18245 10557 18279 10591
rect 13921 10489 13955 10523
rect 1409 10421 1443 10455
rect 2421 10421 2455 10455
rect 5089 10421 5123 10455
rect 5457 10421 5491 10455
rect 6377 10421 6411 10455
rect 7021 10421 7055 10455
rect 7849 10421 7883 10455
rect 10149 10421 10183 10455
rect 10977 10421 11011 10455
rect 12265 10421 12299 10455
rect 12633 10421 12667 10455
rect 14013 10421 14047 10455
rect 14841 10421 14875 10455
rect 17877 10421 17911 10455
rect 2605 10217 2639 10251
rect 3065 10217 3099 10251
rect 3893 10217 3927 10251
rect 8033 10217 8067 10251
rect 18337 10217 18371 10251
rect 2421 10149 2455 10183
rect 4721 10149 4755 10183
rect 13093 10149 13127 10183
rect 17785 10149 17819 10183
rect 3525 10081 3559 10115
rect 4353 10081 4387 10115
rect 4537 10081 4571 10115
rect 5181 10081 5215 10115
rect 5273 10081 5307 10115
rect 6009 10081 6043 10115
rect 6193 10081 6227 10115
rect 6837 10081 6871 10115
rect 6929 10081 6963 10115
rect 7297 10081 7331 10115
rect 8585 10081 8619 10115
rect 8953 10081 8987 10115
rect 11161 10081 11195 10115
rect 12817 10081 12851 10115
rect 13645 10081 13679 10115
rect 14749 10081 14783 10115
rect 15485 10081 15519 10115
rect 16313 10081 16347 10115
rect 17233 10081 17267 10115
rect 1501 10013 1535 10047
rect 1869 10013 1903 10047
rect 2053 10013 2087 10047
rect 2789 10013 2823 10047
rect 5089 10013 5123 10047
rect 7573 10013 7607 10047
rect 8493 10013 8527 10047
rect 9229 10013 9263 10047
rect 11345 10013 11379 10047
rect 11621 10013 11655 10047
rect 13461 10013 13495 10047
rect 14473 10013 14507 10047
rect 16221 10013 16255 10047
rect 17601 10013 17635 10047
rect 18061 10013 18095 10047
rect 2237 9945 2271 9979
rect 3341 9945 3375 9979
rect 4261 9945 4295 9979
rect 10885 9945 10919 9979
rect 12633 9945 12667 9979
rect 18429 9945 18463 9979
rect 1593 9877 1627 9911
rect 3157 9877 3191 9911
rect 5549 9877 5583 9911
rect 5917 9877 5951 9911
rect 6377 9877 6411 9911
rect 6745 9877 6779 9911
rect 7481 9877 7515 9911
rect 7941 9877 7975 9911
rect 8401 9877 8435 9911
rect 10517 9877 10551 9911
rect 10977 9877 11011 9911
rect 12265 9877 12299 9911
rect 12725 9877 12759 9911
rect 13553 9877 13587 9911
rect 14105 9877 14139 9911
rect 14565 9877 14599 9911
rect 14933 9877 14967 9911
rect 15301 9877 15335 9911
rect 15393 9877 15427 9911
rect 15761 9877 15795 9911
rect 16129 9877 16163 9911
rect 16681 9877 16715 9911
rect 17049 9877 17083 9911
rect 17141 9877 17175 9911
rect 17877 9877 17911 9911
rect 2237 9673 2271 9707
rect 5641 9673 5675 9707
rect 6837 9673 6871 9707
rect 8493 9673 8527 9707
rect 9321 9673 9355 9707
rect 10057 9673 10091 9707
rect 10425 9673 10459 9707
rect 11989 9673 12023 9707
rect 13185 9673 13219 9707
rect 14749 9673 14783 9707
rect 15209 9673 15243 9707
rect 16405 9673 16439 9707
rect 18429 9673 18463 9707
rect 1685 9605 1719 9639
rect 3525 9605 3559 9639
rect 5549 9605 5583 9639
rect 6745 9605 6779 9639
rect 14289 9605 14323 9639
rect 14381 9605 14415 9639
rect 15301 9605 15335 9639
rect 15945 9605 15979 9639
rect 16037 9605 16071 9639
rect 16957 9605 16991 9639
rect 1501 9537 1535 9571
rect 2881 9537 2915 9571
rect 4353 9537 4387 9571
rect 7573 9537 7607 9571
rect 8401 9537 8435 9571
rect 9229 9537 9263 9571
rect 11897 9537 11931 9571
rect 12725 9537 12759 9571
rect 13553 9537 13587 9571
rect 16865 9537 16899 9571
rect 17509 9537 17543 9571
rect 18337 9537 18371 9571
rect 1961 9469 1995 9503
rect 2145 9469 2179 9503
rect 3617 9469 3651 9503
rect 3801 9469 3835 9503
rect 4445 9469 4479 9503
rect 4537 9469 4571 9503
rect 4813 9469 4847 9503
rect 5733 9469 5767 9503
rect 6929 9469 6963 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 8677 9469 8711 9503
rect 9413 9469 9447 9503
rect 9781 9469 9815 9503
rect 9965 9469 9999 9503
rect 10517 9469 10551 9503
rect 10793 9469 10827 9503
rect 12081 9469 12115 9503
rect 12817 9469 12851 9503
rect 13001 9469 13035 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 14197 9469 14231 9503
rect 15393 9469 15427 9503
rect 15761 9469 15795 9503
rect 17233 9469 17267 9503
rect 2605 9401 2639 9435
rect 3157 9401 3191 9435
rect 3985 9401 4019 9435
rect 6101 9401 6135 9435
rect 6377 9401 6411 9435
rect 7941 9401 7975 9435
rect 8861 9401 8895 9435
rect 12357 9401 12391 9435
rect 16681 9401 16715 9435
rect 18153 9401 18187 9435
rect 2697 9333 2731 9367
rect 3065 9333 3099 9367
rect 5181 9333 5215 9367
rect 8033 9333 8067 9367
rect 11529 9333 11563 9367
rect 14841 9333 14875 9367
rect 1961 9129 1995 9163
rect 8033 9129 8067 9163
rect 8953 9129 8987 9163
rect 10885 9129 10919 9163
rect 15393 9129 15427 9163
rect 1685 9061 1719 9095
rect 6193 9061 6227 9095
rect 7941 9061 7975 9095
rect 14473 9061 14507 9095
rect 2605 8993 2639 9027
rect 4445 8993 4479 9027
rect 5181 8993 5215 9027
rect 5641 8993 5675 9027
rect 8677 8993 8711 9027
rect 9505 8993 9539 9027
rect 9873 8993 9907 9027
rect 10701 8993 10735 9027
rect 11345 8993 11379 9027
rect 11529 8993 11563 9027
rect 12265 8993 12299 9027
rect 13185 8993 13219 9027
rect 14197 8993 14231 9027
rect 14657 8993 14691 9027
rect 14841 8993 14875 9027
rect 15945 8993 15979 9027
rect 16865 8993 16899 9027
rect 17601 8993 17635 9027
rect 2789 8925 2823 8959
rect 3249 8925 3283 8959
rect 4997 8925 5031 8959
rect 5825 8925 5859 8959
rect 6561 8925 6595 8959
rect 9413 8925 9447 8959
rect 10517 8925 10551 8959
rect 13645 8925 13679 8959
rect 13921 8925 13955 8959
rect 14289 8925 14323 8959
rect 16589 8925 16623 8959
rect 18061 8925 18095 8959
rect 18245 8925 18279 8959
rect 1501 8857 1535 8891
rect 3525 8857 3559 8891
rect 4169 8857 4203 8891
rect 6828 8857 6862 8891
rect 8493 8857 8527 8891
rect 9321 8857 9355 8891
rect 11253 8857 11287 8891
rect 15853 8857 15887 8891
rect 17417 8857 17451 8891
rect 1777 8789 1811 8823
rect 2329 8789 2363 8823
rect 2421 8789 2455 8823
rect 2973 8789 3007 8823
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 4629 8789 4663 8823
rect 5089 8789 5123 8823
rect 5733 8789 5767 8823
rect 6285 8789 6319 8823
rect 8401 8789 8435 8823
rect 10057 8789 10091 8823
rect 10425 8789 10459 8823
rect 13001 8789 13035 8823
rect 13553 8789 13587 8823
rect 14933 8789 14967 8823
rect 15301 8789 15335 8823
rect 15761 8789 15795 8823
rect 16221 8789 16255 8823
rect 16681 8789 16715 8823
rect 17049 8789 17083 8823
rect 17509 8789 17543 8823
rect 17877 8789 17911 8823
rect 18429 8789 18463 8823
rect 1593 8585 1627 8619
rect 2053 8585 2087 8619
rect 2421 8585 2455 8619
rect 3249 8585 3283 8619
rect 3341 8585 3375 8619
rect 4445 8585 4479 8619
rect 6193 8585 6227 8619
rect 8585 8585 8619 8619
rect 10517 8585 10551 8619
rect 13369 8585 13403 8619
rect 14841 8585 14875 8619
rect 16405 8585 16439 8619
rect 16681 8585 16715 8619
rect 17509 8585 17543 8619
rect 17969 8585 18003 8619
rect 1501 8517 1535 8551
rect 3893 8517 3927 8551
rect 15200 8517 15234 8551
rect 17877 8517 17911 8551
rect 1777 8449 1811 8483
rect 2513 8449 2547 8483
rect 4353 8449 4387 8483
rect 4813 8449 4847 8483
rect 5080 8449 5114 8483
rect 6745 8449 6779 8483
rect 7205 8449 7239 8483
rect 7472 8449 7506 8483
rect 9137 8449 9171 8483
rect 9393 8449 9427 8483
rect 11621 8449 11655 8483
rect 11888 8449 11922 8483
rect 13461 8449 13495 8483
rect 13728 8449 13762 8483
rect 14933 8449 14967 8483
rect 17049 8449 17083 8483
rect 17141 8449 17175 8483
rect 18521 8449 18555 8483
rect 2697 8381 2731 8415
rect 3433 8381 3467 8415
rect 4537 8381 4571 8415
rect 6837 8381 6871 8415
rect 6929 8381 6963 8415
rect 17233 8381 17267 8415
rect 18061 8381 18095 8415
rect 1961 8313 1995 8347
rect 3985 8313 4019 8347
rect 6377 8313 6411 8347
rect 8769 8313 8803 8347
rect 13001 8313 13035 8347
rect 13185 8313 13219 8347
rect 16313 8313 16347 8347
rect 18337 8313 18371 8347
rect 2881 8245 2915 8279
rect 8953 8245 8987 8279
rect 1501 8041 1535 8075
rect 2973 8041 3007 8075
rect 4721 8041 4755 8075
rect 5549 8041 5583 8075
rect 7297 8041 7331 8075
rect 9597 8041 9631 8075
rect 17049 8041 17083 8075
rect 18429 8041 18463 8075
rect 2421 7973 2455 8007
rect 12725 7973 12759 8007
rect 16957 7973 16991 8007
rect 3801 7905 3835 7939
rect 4077 7905 4111 7939
rect 4997 7905 5031 7939
rect 5089 7905 5123 7939
rect 10977 7905 11011 7939
rect 11345 7905 11379 7939
rect 17601 7905 17635 7939
rect 1685 7837 1719 7871
rect 2053 7837 2087 7871
rect 2329 7837 2363 7871
rect 2605 7837 2639 7871
rect 3617 7837 3651 7871
rect 4353 7837 4387 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 8769 7837 8803 7871
rect 11601 7837 11635 7871
rect 13645 7837 13679 7871
rect 15485 7837 15519 7871
rect 15577 7837 15611 7871
rect 17417 7837 17451 7871
rect 17877 7837 17911 7871
rect 18245 7837 18279 7871
rect 2789 7769 2823 7803
rect 3341 7769 3375 7803
rect 4261 7769 4295 7803
rect 5181 7769 5215 7803
rect 6184 7769 6218 7803
rect 8524 7769 8558 7803
rect 10732 7769 10766 7803
rect 13921 7769 13955 7803
rect 15218 7769 15252 7803
rect 15844 7769 15878 7803
rect 1869 7701 1903 7735
rect 2145 7701 2179 7735
rect 3065 7701 3099 7735
rect 3433 7701 3467 7735
rect 7389 7701 7423 7735
rect 11161 7701 11195 7735
rect 14105 7701 14139 7735
rect 17509 7701 17543 7735
rect 18061 7701 18095 7735
rect 2973 7497 3007 7531
rect 3341 7497 3375 7531
rect 5089 7497 5123 7531
rect 7941 7497 7975 7531
rect 12909 7497 12943 7531
rect 13737 7497 13771 7531
rect 15393 7497 15427 7531
rect 16221 7497 16255 7531
rect 16681 7497 16715 7531
rect 17049 7497 17083 7531
rect 17141 7497 17175 7531
rect 17969 7497 18003 7531
rect 18337 7497 18371 7531
rect 2053 7429 2087 7463
rect 4445 7429 4479 7463
rect 4997 7429 5031 7463
rect 13093 7429 13127 7463
rect 1685 7361 1719 7395
rect 2145 7361 2179 7395
rect 3801 7361 3835 7395
rect 4353 7361 4387 7395
rect 5549 7361 5583 7395
rect 6828 7361 6862 7395
rect 9137 7361 9171 7395
rect 9404 7361 9438 7395
rect 11529 7361 11563 7395
rect 11785 7361 11819 7395
rect 14850 7361 14884 7395
rect 15117 7361 15151 7395
rect 15209 7361 15243 7395
rect 15485 7361 15519 7395
rect 16129 7361 16163 7395
rect 17877 7361 17911 7395
rect 18521 7361 18555 7395
rect 1961 7293 1995 7327
rect 2697 7293 2731 7327
rect 2881 7293 2915 7327
rect 3893 7293 3927 7327
rect 3985 7293 4019 7327
rect 5181 7293 5215 7327
rect 6561 7293 6595 7327
rect 13277 7293 13311 7327
rect 13461 7293 13495 7327
rect 16313 7293 16347 7327
rect 17325 7293 17359 7327
rect 18061 7293 18095 7327
rect 1501 7225 1535 7259
rect 3433 7225 3467 7259
rect 10517 7225 10551 7259
rect 2513 7157 2547 7191
rect 4629 7157 4663 7191
rect 13645 7157 13679 7191
rect 15669 7157 15703 7191
rect 15761 7157 15795 7191
rect 17509 7157 17543 7191
rect 2605 6953 2639 6987
rect 7297 6953 7331 6987
rect 9965 6953 9999 6987
rect 11437 6953 11471 6987
rect 18429 6953 18463 6987
rect 1501 6885 1535 6919
rect 2237 6885 2271 6919
rect 13369 6885 13403 6919
rect 2329 6817 2363 6851
rect 2973 6817 3007 6851
rect 8769 6817 8803 6851
rect 11345 6817 11379 6851
rect 13001 6817 13035 6851
rect 15485 6817 15519 6851
rect 15577 6817 15611 6851
rect 17601 6817 17635 6851
rect 1685 6749 1719 6783
rect 2053 6749 2087 6783
rect 2789 6749 2823 6783
rect 3985 6749 4019 6783
rect 4445 6749 4479 6783
rect 5917 6749 5951 6783
rect 8513 6749 8547 6783
rect 11078 6749 11112 6783
rect 12817 6749 12851 6783
rect 13461 6749 13495 6783
rect 13737 6749 13771 6783
rect 15229 6749 15263 6783
rect 17509 6749 17543 6783
rect 17877 6749 17911 6783
rect 18245 6749 18279 6783
rect 3157 6681 3191 6715
rect 4261 6681 4295 6715
rect 4712 6681 4746 6715
rect 6184 6681 6218 6715
rect 12550 6681 12584 6715
rect 15822 6681 15856 6715
rect 17417 6681 17451 6715
rect 1869 6613 1903 6647
rect 3249 6613 3283 6647
rect 3617 6613 3651 6647
rect 3801 6613 3835 6647
rect 4077 6613 4111 6647
rect 5825 6613 5859 6647
rect 7389 6613 7423 6647
rect 13185 6613 13219 6647
rect 13645 6613 13679 6647
rect 13921 6613 13955 6647
rect 14105 6613 14139 6647
rect 16957 6613 16991 6647
rect 17049 6613 17083 6647
rect 18061 6613 18095 6647
rect 1777 6409 1811 6443
rect 2789 6409 2823 6443
rect 3249 6409 3283 6443
rect 3985 6409 4019 6443
rect 12449 6409 12483 6443
rect 13461 6409 13495 6443
rect 16313 6409 16347 6443
rect 16865 6409 16899 6443
rect 18429 6409 18463 6443
rect 4077 6341 4111 6375
rect 14596 6341 14630 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2237 6273 2271 6307
rect 2513 6273 2547 6307
rect 3157 6273 3191 6307
rect 4813 6273 4847 6307
rect 5080 6273 5114 6307
rect 7369 6273 7403 6307
rect 9496 6273 9530 6307
rect 11989 6273 12023 6307
rect 12633 6273 12667 6307
rect 13093 6273 13127 6307
rect 13185 6273 13219 6307
rect 14841 6273 14875 6307
rect 14933 6273 14967 6307
rect 15200 6273 15234 6307
rect 16497 6273 16531 6307
rect 16681 6273 16715 6307
rect 17233 6273 17267 6307
rect 17693 6273 17727 6307
rect 17785 6273 17819 6307
rect 18245 6273 18279 6307
rect 3433 6205 3467 6239
rect 3893 6205 3927 6239
rect 6469 6205 6503 6239
rect 7113 6205 7147 6239
rect 9229 6205 9263 6239
rect 12173 6205 12207 6239
rect 17877 6205 17911 6239
rect 2697 6137 2731 6171
rect 11345 6137 11379 6171
rect 13369 6137 13403 6171
rect 1501 6069 1535 6103
rect 2053 6069 2087 6103
rect 2329 6069 2363 6103
rect 4445 6069 4479 6103
rect 4629 6069 4663 6103
rect 6193 6069 6227 6103
rect 6561 6069 6595 6103
rect 6745 6069 6779 6103
rect 6929 6069 6963 6103
rect 8493 6069 8527 6103
rect 10609 6069 10643 6103
rect 11529 6069 11563 6103
rect 11713 6069 11747 6103
rect 12725 6069 12759 6103
rect 12909 6069 12943 6103
rect 17049 6069 17083 6103
rect 17325 6069 17359 6103
rect 2789 5865 2823 5899
rect 4261 5865 4295 5899
rect 11989 5865 12023 5899
rect 13553 5865 13587 5899
rect 15577 5865 15611 5899
rect 3617 5797 3651 5831
rect 6101 5797 6135 5831
rect 12081 5797 12115 5831
rect 2145 5729 2179 5763
rect 2329 5729 2363 5763
rect 3065 5729 3099 5763
rect 4997 5729 5031 5763
rect 5181 5729 5215 5763
rect 5825 5729 5859 5763
rect 13461 5729 13495 5763
rect 16681 5729 16715 5763
rect 17509 5729 17543 5763
rect 18337 5729 18371 5763
rect 1409 5661 1443 5695
rect 1961 5661 1995 5695
rect 2421 5661 2455 5695
rect 3985 5677 4019 5711
rect 4077 5637 4111 5671
rect 5549 5661 5583 5695
rect 7481 5661 7515 5695
rect 9137 5661 9171 5695
rect 9404 5661 9438 5695
rect 10609 5661 10643 5695
rect 13737 5661 13771 5695
rect 14105 5661 14139 5695
rect 15761 5661 15795 5695
rect 16497 5661 16531 5695
rect 3249 5593 3283 5627
rect 4353 5593 4387 5627
rect 7214 5593 7248 5627
rect 10854 5593 10888 5627
rect 13194 5593 13228 5627
rect 14372 5593 14406 5627
rect 16589 5593 16623 5627
rect 1593 5525 1627 5559
rect 1777 5525 1811 5559
rect 3157 5525 3191 5559
rect 3801 5525 3835 5559
rect 4537 5525 4571 5559
rect 4905 5525 4939 5559
rect 5365 5525 5399 5559
rect 5733 5525 5767 5559
rect 10517 5525 10551 5559
rect 13921 5525 13955 5559
rect 15485 5525 15519 5559
rect 15945 5525 15979 5559
rect 16129 5525 16163 5559
rect 16957 5525 16991 5559
rect 17325 5525 17359 5559
rect 17417 5525 17451 5559
rect 17785 5525 17819 5559
rect 18153 5525 18187 5559
rect 18245 5525 18279 5559
rect 1501 5321 1535 5355
rect 3157 5321 3191 5355
rect 3985 5321 4019 5355
rect 4077 5321 4111 5355
rect 4445 5321 4479 5355
rect 4813 5321 4847 5355
rect 4905 5321 4939 5355
rect 5273 5321 5307 5355
rect 8033 5321 8067 5355
rect 9505 5321 9539 5355
rect 15853 5321 15887 5355
rect 17417 5321 17451 5355
rect 18245 5321 18279 5355
rect 18337 5321 18371 5355
rect 5641 5253 5675 5287
rect 6898 5253 6932 5287
rect 17785 5253 17819 5287
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 2329 5185 2363 5219
rect 2605 5185 2639 5219
rect 6653 5185 6687 5219
rect 8125 5185 8159 5219
rect 8381 5185 8415 5219
rect 9965 5185 9999 5219
rect 10232 5185 10266 5219
rect 12642 5185 12676 5219
rect 12909 5185 12943 5219
rect 14114 5185 14148 5219
rect 14381 5185 14415 5219
rect 14473 5185 14507 5219
rect 14740 5185 14774 5219
rect 15945 5185 15979 5219
rect 16497 5185 16531 5219
rect 17049 5185 17083 5219
rect 17877 5185 17911 5219
rect 3249 5117 3283 5151
rect 3341 5117 3375 5151
rect 4261 5117 4295 5151
rect 5089 5117 5123 5151
rect 5733 5117 5767 5151
rect 5825 5117 5859 5151
rect 16773 5117 16807 5151
rect 16957 5117 16991 5151
rect 17601 5117 17635 5151
rect 2421 5049 2455 5083
rect 6193 5049 6227 5083
rect 11529 5049 11563 5083
rect 16129 5049 16163 5083
rect 1869 4981 1903 5015
rect 2145 4981 2179 5015
rect 2789 4981 2823 5015
rect 3617 4981 3651 5015
rect 6377 4981 6411 5015
rect 11345 4981 11379 5015
rect 13001 4981 13035 5015
rect 16313 4981 16347 5015
rect 2881 4777 2915 4811
rect 5825 4777 5859 4811
rect 9045 4777 9079 4811
rect 17969 4777 18003 4811
rect 18429 4777 18463 4811
rect 1777 4709 1811 4743
rect 14105 4709 14139 4743
rect 2237 4641 2271 4675
rect 2329 4641 2363 4675
rect 3341 4641 3375 4675
rect 3525 4641 3559 4675
rect 7205 4641 7239 4675
rect 7389 4641 7423 4675
rect 10425 4641 10459 4675
rect 11345 4641 11379 4675
rect 11713 4641 11747 4675
rect 15485 4641 15519 4675
rect 15669 4641 15703 4675
rect 15853 4641 15887 4675
rect 16957 4641 16991 4675
rect 17325 4641 17359 4675
rect 17509 4641 17543 4675
rect 18153 4641 18187 4675
rect 1685 4573 1719 4607
rect 1961 4573 1995 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 5466 4573 5500 4607
rect 5733 4573 5767 4607
rect 6938 4573 6972 4607
rect 10158 4573 10192 4607
rect 10609 4573 10643 4607
rect 13277 4573 13311 4607
rect 13645 4573 13679 4607
rect 15945 4573 15979 4607
rect 17601 4573 17635 4607
rect 18245 4573 18279 4607
rect 7634 4505 7668 4539
rect 11980 4505 12014 4539
rect 15240 4505 15274 4539
rect 16773 4505 16807 4539
rect 1501 4437 1535 4471
rect 2421 4437 2455 4471
rect 2789 4437 2823 4471
rect 3801 4437 3835 4471
rect 4077 4437 4111 4471
rect 4353 4437 4387 4471
rect 8769 4437 8803 4471
rect 13093 4437 13127 4471
rect 13461 4437 13495 4471
rect 13829 4437 13863 4471
rect 16313 4437 16347 4471
rect 16405 4437 16439 4471
rect 16865 4437 16899 4471
rect 3525 4233 3559 4267
rect 4353 4233 4387 4267
rect 4721 4233 4755 4267
rect 6193 4233 6227 4267
rect 11805 4233 11839 4267
rect 12081 4233 12115 4267
rect 15853 4233 15887 4267
rect 17141 4233 17175 4267
rect 18429 4233 18463 4267
rect 3433 4165 3467 4199
rect 4261 4165 4295 4199
rect 15945 4165 15979 4199
rect 17601 4165 17635 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 3065 4097 3099 4131
rect 5080 4097 5114 4131
rect 6377 4097 6411 4131
rect 7869 4097 7903 4131
rect 8125 4097 8159 4131
rect 9514 4097 9548 4131
rect 9781 4097 9815 4131
rect 9873 4097 9907 4131
rect 10129 4097 10163 4131
rect 11621 4097 11655 4131
rect 11897 4097 11931 4131
rect 12173 4097 12207 4131
rect 12449 4097 12483 4131
rect 12716 4097 12750 4131
rect 14105 4097 14139 4131
rect 14361 4097 14395 4131
rect 17049 4097 17083 4131
rect 17509 4097 17543 4131
rect 18153 4097 18187 4131
rect 18245 4097 18279 4131
rect 2789 4029 2823 4063
rect 3341 4029 3375 4063
rect 4169 4029 4203 4063
rect 4813 4029 4847 4063
rect 15669 4029 15703 4063
rect 16405 4029 16439 4063
rect 17693 4029 17727 4063
rect 1501 3961 1535 3995
rect 6745 3961 6779 3995
rect 8401 3961 8435 3995
rect 15485 3961 15519 3995
rect 16865 3961 16899 3995
rect 17969 3961 18003 3995
rect 1869 3893 1903 3927
rect 2145 3893 2179 3927
rect 2421 3893 2455 3927
rect 2881 3893 2915 3927
rect 3893 3893 3927 3927
rect 6561 3893 6595 3927
rect 8309 3893 8343 3927
rect 11253 3893 11287 3927
rect 12357 3893 12391 3927
rect 13829 3893 13863 3927
rect 14013 3893 14047 3927
rect 16313 3893 16347 3927
rect 3617 3689 3651 3723
rect 6653 3689 6687 3723
rect 12173 3689 12207 3723
rect 16957 3689 16991 3723
rect 17233 3689 17267 3723
rect 17509 3689 17543 3723
rect 18337 3689 18371 3723
rect 2789 3621 2823 3655
rect 6561 3621 6595 3655
rect 9965 3621 9999 3655
rect 11713 3621 11747 3655
rect 3065 3553 3099 3587
rect 4537 3553 4571 3587
rect 8033 3553 8067 3587
rect 11345 3553 11379 3587
rect 13553 3553 13587 3587
rect 15485 3553 15519 3587
rect 15577 3553 15611 3587
rect 17969 3553 18003 3587
rect 18061 3553 18095 3587
rect 1685 3485 1719 3519
rect 1777 3485 1811 3519
rect 2145 3485 2179 3519
rect 2605 3485 2639 3519
rect 3157 3485 3191 3519
rect 3249 3485 3283 3519
rect 3893 3485 3927 3519
rect 4813 3485 4847 3519
rect 5181 3485 5215 3519
rect 7777 3485 7811 3519
rect 8394 3485 8428 3519
rect 8677 3485 8711 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 9597 3485 9631 3519
rect 11529 3485 11563 3519
rect 12081 3485 12115 3519
rect 13286 3485 13320 3519
rect 13921 3485 13955 3519
rect 17417 3485 17451 3519
rect 18521 3485 18555 3519
rect 4445 3417 4479 3451
rect 5426 3417 5460 3451
rect 11100 3417 11134 3451
rect 15240 3417 15274 3451
rect 15822 3417 15856 3451
rect 17877 3417 17911 3451
rect 1501 3349 1535 3383
rect 1961 3349 1995 3383
rect 2329 3349 2363 3383
rect 3985 3349 4019 3383
rect 4353 3349 4387 3383
rect 4997 3349 5031 3383
rect 8217 3349 8251 3383
rect 8493 3349 8527 3383
rect 8953 3349 8987 3383
rect 9229 3349 9263 3383
rect 9781 3349 9815 3383
rect 11897 3349 11931 3383
rect 13737 3349 13771 3383
rect 14105 3349 14139 3383
rect 2973 3145 3007 3179
rect 3893 3145 3927 3179
rect 4261 3145 4295 3179
rect 4813 3145 4847 3179
rect 11989 3145 12023 3179
rect 13461 3145 13495 3179
rect 16313 3145 16347 3179
rect 16957 3145 16991 3179
rect 17325 3145 17359 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 18153 3145 18187 3179
rect 1869 3077 1903 3111
rect 13124 3077 13158 3111
rect 14596 3077 14630 3111
rect 1593 3009 1627 3043
rect 2145 3009 2179 3043
rect 2513 3009 2547 3043
rect 2881 3009 2915 3043
rect 3157 3009 3191 3043
rect 3433 3009 3467 3043
rect 3709 3009 3743 3043
rect 4353 3009 4387 3043
rect 5937 3009 5971 3043
rect 7593 3009 7627 3043
rect 7849 3009 7883 3043
rect 8401 3009 8435 3043
rect 8749 3009 8783 3043
rect 9965 3009 9999 3043
rect 10232 3009 10266 3043
rect 11529 3009 11563 3043
rect 13369 3009 13403 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 15200 3009 15234 3043
rect 16865 3009 16899 3043
rect 18245 3009 18279 3043
rect 4169 2941 4203 2975
rect 6193 2941 6227 2975
rect 8033 2941 8067 2975
rect 8493 2941 8527 2975
rect 17509 2941 17543 2975
rect 18337 2941 18371 2975
rect 3341 2873 3375 2907
rect 11713 2873 11747 2907
rect 16497 2873 16531 2907
rect 1409 2805 1443 2839
rect 2329 2805 2363 2839
rect 2697 2805 2731 2839
rect 3617 2805 3651 2839
rect 4721 2805 4755 2839
rect 6469 2805 6503 2839
rect 8217 2805 8251 2839
rect 9873 2805 9907 2839
rect 11345 2805 11379 2839
rect 16681 2805 16715 2839
rect 1593 2601 1627 2635
rect 3893 2601 3927 2635
rect 4169 2601 4203 2635
rect 5917 2601 5951 2635
rect 9137 2601 9171 2635
rect 11529 2601 11563 2635
rect 13553 2601 13587 2635
rect 16037 2601 16071 2635
rect 16313 2601 16347 2635
rect 17233 2601 17267 2635
rect 18061 2601 18095 2635
rect 18429 2601 18463 2635
rect 2605 2533 2639 2567
rect 6193 2533 6227 2567
rect 8585 2533 8619 2567
rect 13185 2533 13219 2567
rect 15761 2533 15795 2567
rect 4537 2465 4571 2499
rect 4629 2465 4663 2499
rect 5365 2465 5399 2499
rect 5457 2465 5491 2499
rect 9597 2465 9631 2499
rect 9781 2465 9815 2499
rect 11345 2465 11379 2499
rect 12909 2465 12943 2499
rect 15485 2465 15519 2499
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 2421 2397 2455 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 8401 2397 8435 2431
rect 8769 2397 8803 2431
rect 9045 2397 9079 2431
rect 13001 2397 13035 2431
rect 13369 2397 13403 2431
rect 13737 2397 13771 2431
rect 15577 2397 15611 2431
rect 16221 2397 16255 2431
rect 16497 2397 16531 2431
rect 16773 2397 16807 2431
rect 17417 2397 17451 2431
rect 17509 2397 17543 2431
rect 17877 2397 17911 2431
rect 18245 2397 18279 2431
rect 5549 2329 5583 2363
rect 8156 2329 8190 2363
rect 9505 2329 9539 2363
rect 11078 2329 11112 2363
rect 12642 2329 12676 2363
rect 15218 2329 15252 2363
rect 1869 2261 1903 2295
rect 2237 2261 2271 2295
rect 3065 2261 3099 2295
rect 3525 2261 3559 2295
rect 5089 2261 5123 2295
rect 6561 2261 6595 2295
rect 6837 2261 6871 2295
rect 7021 2261 7055 2295
rect 9965 2261 9999 2295
rect 13921 2261 13955 2295
rect 14105 2261 14139 2295
rect 16957 2261 16991 2295
rect 17693 2261 17727 2295
<< metal1 >>
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 6546 15008 6552 15020
rect 2372 14980 6552 15008
rect 2372 14968 2378 14980
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 15286 14940 15292 14952
rect 5960 14912 15292 14940
rect 5960 14900 5966 14912
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 3602 14832 3608 14884
rect 3660 14872 3666 14884
rect 6914 14872 6920 14884
rect 3660 14844 6920 14872
rect 3660 14832 3666 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 5442 14804 5448 14816
rect 4488 14776 5448 14804
rect 4488 14764 4494 14776
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 16206 14804 16212 14816
rect 15252 14776 16212 14804
rect 15252 14764 15258 14776
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 5718 14600 5724 14612
rect 2832 14572 5396 14600
rect 5679 14572 5724 14600
rect 2832 14560 2838 14572
rect 2240 14504 5304 14532
rect 2240 14476 2268 14504
rect 2222 14464 2228 14476
rect 2135 14436 2228 14464
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 3145 14467 3203 14473
rect 3145 14464 3157 14467
rect 2832 14436 3157 14464
rect 2832 14424 2838 14436
rect 3145 14433 3157 14436
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 3510 14424 3516 14476
rect 3568 14464 3574 14476
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 3568 14436 5181 14464
rect 3568 14424 3574 14436
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 2884 14260 2912 14359
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 4062 14396 4068 14408
rect 3016 14368 4068 14396
rect 3016 14356 3022 14368
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4246 14356 4252 14408
rect 4304 14396 4310 14408
rect 4341 14399 4399 14405
rect 4341 14396 4353 14399
rect 4304 14368 4353 14396
rect 4304 14356 4310 14368
rect 4341 14365 4353 14368
rect 4387 14365 4399 14399
rect 4341 14359 4399 14365
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 4724 14405 4752 14436
rect 5169 14433 5181 14436
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4488 14368 4629 14396
rect 4488 14356 4494 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 5276 14396 5304 14504
rect 5368 14464 5396 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6546 14600 6552 14612
rect 6507 14572 6552 14600
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7524 14572 7665 14600
rect 7524 14560 7530 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 10134 14600 10140 14612
rect 10095 14572 10140 14600
rect 7653 14563 7711 14569
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 6917 14535 6975 14541
rect 6917 14532 6929 14535
rect 5592 14504 6929 14532
rect 5592 14492 5598 14504
rect 6917 14501 6929 14504
rect 6963 14501 6975 14535
rect 6917 14495 6975 14501
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 5368 14436 6745 14464
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 5534 14396 5540 14408
rect 4709 14359 4767 14365
rect 4816 14368 5120 14396
rect 5276 14368 5540 14396
rect 3050 14288 3056 14340
rect 3108 14328 3114 14340
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 3108 14300 3433 14328
rect 3108 14288 3114 14300
rect 3421 14297 3433 14300
rect 3467 14328 3479 14331
rect 4816 14328 4844 14368
rect 3467 14300 4844 14328
rect 5092 14328 5120 14368
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5902 14396 5908 14408
rect 5863 14368 5908 14396
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 7668 14396 7696 14563
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12345 14603 12403 14609
rect 12345 14600 12357 14603
rect 12032 14572 12357 14600
rect 12032 14560 12038 14572
rect 12345 14569 12357 14572
rect 12391 14569 12403 14603
rect 14550 14600 14556 14612
rect 14511 14572 14556 14600
rect 12345 14563 12403 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 15028 14572 16574 14600
rect 14369 14535 14427 14541
rect 14369 14501 14381 14535
rect 14415 14532 14427 14535
rect 15028 14532 15056 14572
rect 14415 14504 15056 14532
rect 15105 14535 15163 14541
rect 14415 14501 14427 14504
rect 14369 14495 14427 14501
rect 15105 14501 15117 14535
rect 15151 14532 15163 14535
rect 15470 14532 15476 14544
rect 15151 14504 15476 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14501 15623 14535
rect 16546 14532 16574 14572
rect 16546 14504 17724 14532
rect 15565 14495 15623 14501
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15194 14464 15200 14476
rect 14967 14436 15200 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15580 14464 15608 14495
rect 15654 14464 15660 14476
rect 15580 14436 15660 14464
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 16850 14464 16856 14476
rect 15764 14436 16856 14464
rect 7837 14399 7895 14405
rect 7837 14396 7849 14399
rect 7668 14368 7849 14396
rect 7837 14365 7849 14368
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10870 14396 10876 14408
rect 10367 14368 10876 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 12802 14396 12808 14408
rect 12575 14368 12808 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14737 14399 14795 14405
rect 14737 14396 14749 14399
rect 13872 14368 14749 14396
rect 13872 14356 13878 14368
rect 14737 14365 14749 14368
rect 14783 14396 14795 14399
rect 15378 14396 15384 14408
rect 14783 14368 15384 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 15764 14405 15792 14436
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 17696 14408 17724 14504
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15519 14368 15761 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 16390 14396 16396 14408
rect 15749 14359 15807 14365
rect 15948 14368 16396 14396
rect 6365 14331 6423 14337
rect 6365 14328 6377 14331
rect 5092 14300 6377 14328
rect 3467 14297 3479 14300
rect 3421 14291 3479 14297
rect 6365 14297 6377 14300
rect 6411 14297 6423 14331
rect 6365 14291 6423 14297
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 15194 14328 15200 14340
rect 8168 14300 15200 14328
rect 8168 14288 8174 14300
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15289 14331 15347 14337
rect 15289 14297 15301 14331
rect 15335 14328 15347 14331
rect 15948 14328 15976 14368
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16546 14368 16773 14396
rect 15335 14300 15976 14328
rect 15335 14297 15347 14300
rect 15289 14291 15347 14297
rect 16022 14288 16028 14340
rect 16080 14328 16086 14340
rect 16080 14300 16125 14328
rect 16080 14288 16086 14300
rect 16206 14288 16212 14340
rect 16264 14328 16270 14340
rect 16546 14328 16574 14368
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 17034 14396 17040 14408
rect 16995 14368 17040 14396
rect 16761 14359 16819 14365
rect 17034 14356 17040 14368
rect 17092 14356 17098 14408
rect 17678 14396 17684 14408
rect 17639 14368 17684 14396
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 17957 14399 18015 14405
rect 17957 14396 17969 14399
rect 17920 14368 17969 14396
rect 17920 14356 17926 14368
rect 17957 14365 17969 14368
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 16264 14300 16574 14328
rect 16264 14288 16270 14300
rect 3142 14260 3148 14272
rect 2884 14232 3148 14260
rect 3142 14220 3148 14232
rect 3200 14220 3206 14272
rect 3326 14260 3332 14272
rect 3287 14232 3332 14260
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 4890 14260 4896 14272
rect 4851 14232 4896 14260
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5040 14232 5085 14260
rect 5040 14220 5046 14232
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 5353 14263 5411 14269
rect 5353 14260 5365 14263
rect 5316 14232 5365 14260
rect 5316 14220 5322 14232
rect 5353 14229 5365 14232
rect 5399 14229 5411 14263
rect 5353 14223 5411 14229
rect 5442 14220 5448 14272
rect 5500 14260 5506 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5500 14232 6009 14260
rect 5500 14220 5506 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 5997 14223 6055 14229
rect 8021 14263 8079 14269
rect 8021 14229 8033 14263
rect 8067 14260 8079 14263
rect 10226 14260 10232 14272
rect 8067 14232 10232 14260
rect 8067 14229 8079 14232
rect 8021 14223 8079 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 14148 14232 15945 14260
rect 14148 14220 14154 14232
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 15933 14223 15991 14229
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 16172 14232 16313 14260
rect 16172 14220 16178 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4430 14056 4436 14068
rect 4203 14028 4436 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4571 14028 4997 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 4985 14019 5043 14025
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 5316 14028 5365 14056
rect 5316 14016 5322 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 5353 14019 5411 14025
rect 5445 14059 5503 14065
rect 5445 14025 5457 14059
rect 5491 14056 5503 14059
rect 5994 14056 6000 14068
rect 5491 14028 6000 14056
rect 5491 14025 5503 14028
rect 5445 14019 5503 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6914 14056 6920 14068
rect 6196 14028 6592 14056
rect 6875 14028 6920 14056
rect 6196 13988 6224 14028
rect 2746 13960 6224 13988
rect 6564 13988 6592 14028
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 12802 14056 12808 14068
rect 12763 14028 12808 14056
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 12912 14028 17417 14056
rect 7101 13991 7159 13997
rect 7101 13988 7113 13991
rect 6564 13960 7113 13988
rect 2746 13932 2774 13960
rect 7101 13957 7113 13960
rect 7147 13957 7159 13991
rect 12912 13988 12940 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 7101 13951 7159 13957
rect 9646 13960 12940 13988
rect 13219 13991 13277 13997
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13920 2283 13923
rect 2746 13920 2780 13932
rect 2271 13892 2780 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 2958 13880 2964 13932
rect 3016 13920 3022 13932
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 3016 13892 3341 13920
rect 3016 13880 3022 13892
rect 3329 13889 3341 13892
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3694 13880 3700 13932
rect 3752 13920 3758 13932
rect 3752 13892 3797 13920
rect 3752 13880 3758 13892
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 4120 13892 6377 13920
rect 4120 13880 4126 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 1762 13812 1768 13864
rect 1820 13852 1826 13864
rect 1949 13855 2007 13861
rect 1949 13852 1961 13855
rect 1820 13824 1961 13852
rect 1820 13812 1826 13824
rect 1949 13821 1961 13824
rect 1995 13821 2007 13855
rect 2866 13852 2872 13864
rect 2827 13824 2872 13852
rect 1949 13815 2007 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 3418 13852 3424 13864
rect 3191 13824 3424 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3602 13852 3608 13864
rect 3559 13824 3608 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 3881 13855 3939 13861
rect 3881 13852 3893 13855
rect 3844 13824 3893 13852
rect 3844 13812 3850 13824
rect 3881 13821 3893 13824
rect 3927 13821 3939 13855
rect 4614 13852 4620 13864
rect 4575 13824 4620 13852
rect 3881 13815 3939 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4706 13812 4712 13864
rect 4764 13852 4770 13864
rect 4982 13852 4988 13864
rect 4764 13824 4988 13852
rect 4764 13812 4770 13824
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5132 13824 5641 13852
rect 5132 13812 5138 13824
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5675 13824 5825 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5813 13821 5825 13824
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 8938 13852 8944 13864
rect 6052 13824 8944 13852
rect 6052 13812 6058 13824
rect 8938 13812 8944 13824
rect 8996 13852 9002 13864
rect 9646 13852 9674 13960
rect 13219 13957 13231 13991
rect 13265 13988 13277 13991
rect 15013 13991 15071 13997
rect 15013 13988 15025 13991
rect 13265 13960 15025 13988
rect 13265 13957 13277 13960
rect 13219 13951 13277 13957
rect 15013 13957 15025 13960
rect 15059 13957 15071 13991
rect 15654 13988 15660 14000
rect 15013 13951 15071 13957
rect 15212 13960 15660 13988
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12952 13892 13001 13920
rect 12952 13880 12958 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 13116 13923 13174 13929
rect 13116 13920 13128 13923
rect 12989 13883 13047 13889
rect 13096 13889 13128 13920
rect 13162 13920 13174 13923
rect 13814 13920 13820 13932
rect 13162 13892 13820 13920
rect 13162 13889 13174 13892
rect 13096 13883 13174 13889
rect 8996 13824 9674 13852
rect 10965 13855 11023 13861
rect 8996 13812 9002 13824
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 13096 13852 13124 13883
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 15212 13929 15240 13960
rect 15654 13948 15660 13960
rect 15712 13948 15718 14000
rect 15749 13991 15807 13997
rect 15749 13957 15761 13991
rect 15795 13988 15807 13991
rect 17126 13988 17132 14000
rect 15795 13960 17132 13988
rect 15795 13957 15807 13960
rect 15749 13951 15807 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 17494 13988 17500 14000
rect 17455 13960 17500 13988
rect 17494 13948 17500 13960
rect 17552 13948 17558 14000
rect 15197 13923 15255 13929
rect 15197 13889 15209 13923
rect 15243 13889 15255 13923
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 15197 13883 15255 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15930 13920 15936 13932
rect 15891 13892 15936 13920
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16022 13880 16028 13932
rect 16080 13880 16086 13932
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16298 13920 16304 13932
rect 16163 13892 16304 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16298 13880 16304 13892
rect 16356 13920 16362 13932
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 16356 13892 16405 13920
rect 16356 13880 16362 13892
rect 16393 13889 16405 13892
rect 16439 13889 16451 13923
rect 16666 13920 16672 13932
rect 16627 13892 16672 13920
rect 16393 13883 16451 13889
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 13538 13852 13544 13864
rect 11011 13824 13124 13852
rect 13499 13824 13544 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 16040 13852 16068 13880
rect 14056 13824 16068 13852
rect 16209 13855 16267 13861
rect 14056 13812 14062 13824
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16209 13815 16267 13821
rect 16316 13824 16957 13852
rect 1118 13744 1124 13796
rect 1176 13784 1182 13796
rect 3973 13787 4031 13793
rect 3973 13784 3985 13787
rect 1176 13756 2774 13784
rect 1176 13744 1182 13756
rect 2746 13716 2774 13756
rect 3804 13756 3985 13784
rect 3050 13716 3056 13728
rect 2746 13688 3056 13716
rect 3050 13676 3056 13688
rect 3108 13716 3114 13728
rect 3804 13716 3832 13756
rect 3973 13753 3985 13756
rect 4019 13753 4031 13787
rect 3973 13747 4031 13753
rect 4062 13744 4068 13796
rect 4120 13784 4126 13796
rect 6549 13787 6607 13793
rect 6549 13784 6561 13787
rect 4120 13756 5028 13784
rect 4120 13744 4126 13756
rect 3108 13688 3832 13716
rect 3108 13676 3114 13688
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4890 13716 4896 13728
rect 3936 13688 4896 13716
rect 3936 13676 3942 13688
rect 4890 13676 4896 13688
rect 4948 13676 4954 13728
rect 5000 13716 5028 13756
rect 5644 13756 6561 13784
rect 5644 13716 5672 13756
rect 6549 13753 6561 13756
rect 6595 13753 6607 13787
rect 15286 13784 15292 13796
rect 15247 13756 15292 13784
rect 6549 13747 6607 13753
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 16114 13744 16120 13796
rect 16172 13784 16178 13796
rect 16224 13784 16252 13815
rect 16172 13756 16252 13784
rect 16172 13744 16178 13756
rect 5000 13688 5672 13716
rect 6454 13676 6460 13728
rect 6512 13716 6518 13728
rect 6733 13719 6791 13725
rect 6733 13716 6745 13719
rect 6512 13688 6745 13716
rect 6512 13676 6518 13688
rect 6733 13685 6745 13688
rect 6779 13685 6791 13719
rect 6733 13679 6791 13685
rect 10781 13719 10839 13725
rect 10781 13685 10793 13719
rect 10827 13716 10839 13719
rect 10870 13716 10876 13728
rect 10827 13688 10876 13716
rect 10827 13685 10839 13688
rect 10781 13679 10839 13685
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15654 13716 15660 13728
rect 15252 13688 15660 13716
rect 15252 13676 15258 13688
rect 15654 13676 15660 13688
rect 15712 13716 15718 13728
rect 16316 13716 16344 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 17678 13852 17684 13864
rect 17639 13824 17684 13852
rect 16945 13815 17003 13821
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18322 13852 18328 13864
rect 18003 13824 18328 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 16850 13784 16856 13796
rect 16811 13756 16856 13784
rect 16850 13744 16856 13756
rect 16908 13744 16914 13796
rect 15712 13688 16344 13716
rect 15712 13676 15718 13688
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3418 13512 3424 13524
rect 3108 13484 3424 13512
rect 3108 13472 3114 13484
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 4614 13512 4620 13524
rect 3651 13484 4620 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 6270 13512 6276 13524
rect 4816 13484 6276 13512
rect 4816 13444 4844 13484
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 6822 13512 6828 13524
rect 6783 13484 6828 13512
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 1964 13416 4844 13444
rect 1964 13385 1992 13416
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 17770 13444 17776 13456
rect 16816 13416 17776 13444
rect 16816 13404 16822 13416
rect 17770 13404 17776 13416
rect 17828 13404 17834 13456
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13345 2007 13379
rect 3050 13376 3056 13388
rect 2963 13348 3056 13376
rect 1949 13339 2007 13345
rect 3050 13336 3056 13348
rect 3108 13376 3114 13388
rect 3878 13376 3884 13388
rect 3108 13348 3884 13376
rect 3108 13336 3114 13348
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 5123 13348 5917 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 5905 13345 5917 13348
rect 5951 13345 5963 13379
rect 5905 13339 5963 13345
rect 2222 13308 2228 13320
rect 2183 13280 2228 13308
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 3142 13308 3148 13320
rect 3103 13280 3148 13308
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3418 13268 3424 13320
rect 3476 13308 3482 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3476 13280 3801 13308
rect 3476 13268 3482 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5092 13308 5120 13339
rect 6086 13336 6092 13388
rect 6144 13376 6150 13388
rect 6914 13376 6920 13388
rect 6144 13348 6920 13376
rect 6144 13336 6150 13348
rect 6914 13336 6920 13348
rect 6972 13376 6978 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 6972 13348 7573 13376
rect 6972 13336 6978 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 15013 13379 15071 13385
rect 15013 13345 15025 13379
rect 15059 13376 15071 13379
rect 17954 13376 17960 13388
rect 15059 13348 17724 13376
rect 17915 13348 17960 13376
rect 15059 13345 15071 13348
rect 15013 13339 15071 13345
rect 17696 13320 17724 13348
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 5718 13308 5724 13320
rect 4764 13280 5120 13308
rect 5679 13280 5724 13308
rect 4764 13268 4770 13280
rect 5718 13268 5724 13280
rect 5776 13308 5782 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 5776 13280 6469 13308
rect 5776 13268 5782 13280
rect 6457 13277 6469 13280
rect 6503 13308 6515 13311
rect 6546 13308 6552 13320
rect 6503 13280 6552 13308
rect 6503 13277 6515 13280
rect 6457 13271 6515 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 6880 13280 7389 13308
rect 6880 13268 6886 13280
rect 7377 13277 7389 13280
rect 7423 13308 7435 13311
rect 15102 13308 15108 13320
rect 7423 13280 9674 13308
rect 15063 13280 15108 13308
rect 7423 13277 7435 13280
rect 7377 13271 7435 13277
rect 2409 13243 2467 13249
rect 2409 13209 2421 13243
rect 2455 13240 2467 13243
rect 2866 13240 2872 13252
rect 2455 13212 2872 13240
rect 2455 13209 2467 13212
rect 2409 13203 2467 13209
rect 2866 13200 2872 13212
rect 2924 13240 2930 13252
rect 3694 13240 3700 13252
rect 2924 13212 3700 13240
rect 2924 13200 2930 13212
rect 3694 13200 3700 13212
rect 3752 13200 3758 13252
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 4433 13243 4491 13249
rect 4212 13212 4257 13240
rect 4212 13200 4218 13212
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 4893 13243 4951 13249
rect 4893 13240 4905 13243
rect 4479 13212 4905 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 4893 13209 4905 13212
rect 4939 13209 4951 13243
rect 5810 13240 5816 13252
rect 5771 13212 5816 13240
rect 4893 13203 4951 13209
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 5994 13200 6000 13252
rect 6052 13240 6058 13252
rect 6641 13243 6699 13249
rect 6641 13240 6653 13243
rect 6052 13212 6653 13240
rect 6052 13200 6058 13212
rect 6641 13209 6653 13212
rect 6687 13209 6699 13243
rect 9646 13240 9674 13280
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 17313 13311 17371 13317
rect 17313 13308 17325 13311
rect 16546 13280 17325 13308
rect 13262 13240 13268 13252
rect 9646 13212 13268 13240
rect 6641 13203 6699 13209
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 15289 13243 15347 13249
rect 15289 13209 15301 13243
rect 15335 13240 15347 13243
rect 15378 13240 15384 13252
rect 15335 13212 15384 13240
rect 15335 13209 15347 13212
rect 15289 13203 15347 13209
rect 15378 13200 15384 13212
rect 15436 13200 15442 13252
rect 1210 13132 1216 13184
rect 1268 13172 1274 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 1268 13144 2513 13172
rect 1268 13132 1274 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2501 13135 2559 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 3016 13144 3249 13172
rect 3016 13132 3022 13144
rect 3237 13141 3249 13144
rect 3283 13141 3295 13175
rect 3237 13135 3295 13141
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 4028 13144 4073 13172
rect 4028 13132 4034 13144
rect 4522 13132 4528 13184
rect 4580 13172 4586 13184
rect 4982 13172 4988 13184
rect 4580 13144 4625 13172
rect 4943 13144 4988 13172
rect 4580 13132 4586 13144
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 5353 13175 5411 13181
rect 5353 13172 5365 13175
rect 5132 13144 5365 13172
rect 5132 13132 5138 13144
rect 5353 13141 5365 13144
rect 5399 13141 5411 13175
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 5353 13135 5411 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 7006 13172 7012 13184
rect 6967 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7469 13175 7527 13181
rect 7469 13141 7481 13175
rect 7515 13172 7527 13175
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7515 13144 7941 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7929 13141 7941 13144
rect 7975 13172 7987 13175
rect 11146 13172 11152 13184
rect 7975 13144 11152 13172
rect 7975 13141 7987 13144
rect 7929 13135 7987 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 16546 13172 16574 13280
rect 17313 13277 17325 13280
rect 17359 13277 17371 13311
rect 17678 13308 17684 13320
rect 17639 13280 17684 13308
rect 17313 13271 17371 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 16945 13243 17003 13249
rect 16945 13209 16957 13243
rect 16991 13240 17003 13243
rect 17494 13240 17500 13252
rect 16991 13212 17356 13240
rect 17455 13212 17500 13240
rect 16991 13209 17003 13212
rect 16945 13203 17003 13209
rect 17218 13172 17224 13184
rect 14884 13144 16574 13172
rect 17179 13144 17224 13172
rect 14884 13132 14890 13144
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 17328 13172 17356 13212
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18782 13172 18788 13184
rect 17328 13144 18788 13172
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 2130 12928 2136 12980
rect 2188 12968 2194 12980
rect 3050 12968 3056 12980
rect 2188 12940 3056 12968
rect 2188 12928 2194 12940
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3510 12968 3516 12980
rect 3471 12940 3516 12968
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 3878 12968 3884 12980
rect 3839 12940 3884 12968
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4522 12968 4528 12980
rect 4483 12940 4528 12968
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 4617 12971 4675 12977
rect 4617 12937 4629 12971
rect 4663 12968 4675 12971
rect 5074 12968 5080 12980
rect 4663 12940 5080 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 6181 12971 6239 12977
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6733 12971 6791 12977
rect 6733 12968 6745 12971
rect 6227 12940 6745 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6733 12937 6745 12940
rect 6779 12937 6791 12971
rect 6733 12931 6791 12937
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 7285 12971 7343 12977
rect 7285 12968 7297 12971
rect 6880 12940 7297 12968
rect 6880 12928 6886 12940
rect 7285 12937 7297 12940
rect 7331 12937 7343 12971
rect 7285 12931 7343 12937
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7432 12940 7665 12968
rect 7432 12928 7438 12940
rect 7653 12937 7665 12940
rect 7699 12968 7711 12971
rect 8573 12971 8631 12977
rect 8573 12968 8585 12971
rect 7699 12940 8585 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 8573 12937 8585 12940
rect 8619 12937 8631 12971
rect 8573 12931 8631 12937
rect 15749 12971 15807 12977
rect 15749 12937 15761 12971
rect 15795 12968 15807 12971
rect 17586 12968 17592 12980
rect 15795 12940 17592 12968
rect 15795 12937 15807 12940
rect 15749 12931 15807 12937
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 6454 12900 6460 12912
rect 2240 12872 6460 12900
rect 2240 12776 2268 12872
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 7006 12900 7012 12912
rect 6687 12872 7012 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 8113 12903 8171 12909
rect 8113 12900 8125 12903
rect 7116 12872 8125 12900
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 2556 12804 2697 12832
rect 2556 12792 2562 12804
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 4890 12832 4896 12844
rect 3375 12804 4896 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5626 12832 5632 12844
rect 5399 12804 5632 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 7116 12832 7144 12872
rect 8113 12869 8125 12872
rect 8159 12869 8171 12903
rect 13446 12900 13452 12912
rect 13407 12872 13452 12900
rect 8113 12863 8171 12869
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 16117 12903 16175 12909
rect 16117 12869 16129 12903
rect 16163 12900 16175 12903
rect 17494 12900 17500 12912
rect 16163 12872 17500 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 5859 12804 7144 12832
rect 7745 12835 7803 12841
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 7791 12804 8493 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8481 12801 8493 12804
rect 8527 12832 8539 12835
rect 10594 12832 10600 12844
rect 8527 12804 10600 12832
rect 8527 12801 8539 12804
rect 8481 12795 8539 12801
rect 10594 12792 10600 12804
rect 10652 12832 10658 12844
rect 12618 12832 12624 12844
rect 10652 12804 12624 12832
rect 10652 12792 10658 12804
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12832 13415 12835
rect 13817 12835 13875 12841
rect 13817 12832 13829 12835
rect 13403 12804 13829 12832
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 13817 12801 13829 12804
rect 13863 12801 13875 12835
rect 16298 12832 16304 12844
rect 16259 12804 16304 12832
rect 13817 12795 13875 12801
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17310 12832 17316 12844
rect 16991 12804 17316 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12733 2007 12767
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 1949 12727 2007 12733
rect 1964 12696 1992 12727
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2406 12764 2412 12776
rect 2367 12736 2412 12764
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4580 12736 4721 12764
rect 4580 12724 4586 12736
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 6362 12764 6368 12776
rect 5767 12736 6368 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 2774 12696 2780 12708
rect 1964 12668 2780 12696
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 2958 12656 2964 12708
rect 3016 12696 3022 12708
rect 3145 12699 3203 12705
rect 3145 12696 3157 12699
rect 3016 12668 3157 12696
rect 3016 12656 3022 12668
rect 3145 12665 3157 12668
rect 3191 12665 3203 12699
rect 3970 12696 3976 12708
rect 3145 12659 3203 12665
rect 3344 12668 3976 12696
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3344 12628 3372 12668
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 5552 12696 5580 12727
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 6549 12767 6607 12773
rect 6549 12733 6561 12767
rect 6595 12764 6607 12767
rect 7374 12764 7380 12776
rect 6595 12736 7380 12764
rect 6595 12733 6607 12736
rect 6549 12727 6607 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7524 12736 7849 12764
rect 7524 12724 7530 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 9306 12764 9312 12776
rect 9267 12736 9312 12764
rect 7837 12727 7895 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 14642 12764 14648 12776
rect 13679 12736 14648 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 17678 12764 17684 12776
rect 15979 12736 17684 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 17957 12767 18015 12773
rect 17957 12733 17969 12767
rect 18003 12733 18015 12767
rect 17957 12727 18015 12733
rect 6086 12696 6092 12708
rect 5552 12668 6092 12696
rect 6086 12656 6092 12668
rect 6144 12656 6150 12708
rect 9214 12656 9220 12708
rect 9272 12696 9278 12708
rect 9861 12699 9919 12705
rect 9861 12696 9873 12699
rect 9272 12668 9873 12696
rect 9272 12656 9278 12668
rect 9861 12665 9873 12668
rect 9907 12696 9919 12699
rect 16114 12696 16120 12708
rect 9907 12668 16120 12696
rect 9907 12665 9919 12668
rect 9861 12659 9919 12665
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 17972 12696 18000 12727
rect 16224 12668 18000 12696
rect 3099 12600 3372 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 3697 12631 3755 12637
rect 3697 12628 3709 12631
rect 3568 12600 3709 12628
rect 3568 12588 3574 12600
rect 3697 12597 3709 12600
rect 3743 12597 3755 12631
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 3697 12591 3755 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6730 12628 6736 12640
rect 6052 12600 6736 12628
rect 6052 12588 6058 12600
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 7101 12631 7159 12637
rect 7101 12628 7113 12631
rect 6880 12600 7113 12628
rect 6880 12588 6886 12600
rect 7101 12597 7113 12600
rect 7147 12597 7159 12631
rect 9674 12628 9680 12640
rect 9635 12600 9680 12628
rect 7101 12591 7159 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 16224 12628 16252 12668
rect 13780 12600 16252 12628
rect 13780 12588 13786 12600
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 16448 12600 16493 12628
rect 16448 12588 16454 12600
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 17129 12631 17187 12637
rect 17129 12628 17141 12631
rect 17092 12600 17141 12628
rect 17092 12588 17098 12600
rect 17129 12597 17141 12600
rect 17175 12597 17187 12631
rect 17129 12591 17187 12597
rect 17405 12631 17463 12637
rect 17405 12597 17417 12631
rect 17451 12628 17463 12631
rect 17494 12628 17500 12640
rect 17451 12600 17500 12628
rect 17451 12597 17463 12600
rect 17405 12591 17463 12597
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 17586 12588 17592 12640
rect 17644 12628 17650 12640
rect 18138 12628 18144 12640
rect 17644 12600 18144 12628
rect 17644 12588 17650 12600
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2501 12427 2559 12433
rect 2501 12393 2513 12427
rect 2547 12424 2559 12427
rect 2866 12424 2872 12436
rect 2547 12396 2872 12424
rect 2547 12393 2559 12396
rect 2501 12387 2559 12393
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 5074 12424 5080 12436
rect 4304 12396 5080 12424
rect 4304 12384 4310 12396
rect 5074 12384 5080 12396
rect 5132 12424 5138 12436
rect 9674 12424 9680 12436
rect 5132 12396 9680 12424
rect 5132 12384 5138 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10336 12396 10701 12424
rect 8113 12359 8171 12365
rect 8113 12356 8125 12359
rect 2240 12328 8125 12356
rect 2240 12232 2268 12328
rect 8113 12325 8125 12328
rect 8159 12325 8171 12359
rect 8113 12319 8171 12325
rect 10226 12316 10232 12368
rect 10284 12356 10290 12368
rect 10336 12356 10364 12396
rect 10689 12393 10701 12396
rect 10735 12424 10747 12427
rect 12526 12424 12532 12436
rect 10735 12396 12532 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 13722 12424 13728 12436
rect 13504 12396 13728 12424
rect 13504 12384 13510 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 15013 12427 15071 12433
rect 15013 12393 15025 12427
rect 15059 12424 15071 12427
rect 17862 12424 17868 12436
rect 15059 12396 17868 12424
rect 15059 12393 15071 12396
rect 15013 12387 15071 12393
rect 10284 12328 10364 12356
rect 10284 12316 10290 12328
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 12434 12356 12440 12368
rect 10468 12328 12440 12356
rect 10468 12316 10474 12328
rect 12434 12316 12440 12328
rect 12492 12316 12498 12368
rect 14090 12316 14096 12368
rect 14148 12356 14154 12368
rect 14826 12356 14832 12368
rect 14148 12328 14832 12356
rect 14148 12316 14154 12328
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 3510 12288 3516 12300
rect 3471 12260 3516 12288
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 3752 12260 4353 12288
rect 3752 12248 3758 12260
rect 4341 12257 4353 12260
rect 4387 12288 4399 12291
rect 4522 12288 4528 12300
rect 4387 12260 4528 12288
rect 4387 12257 4399 12260
rect 4341 12251 4399 12257
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12257 4767 12291
rect 4890 12288 4896 12300
rect 4851 12260 4896 12288
rect 4709 12251 4767 12257
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2222 12220 2228 12232
rect 2183 12192 2228 12220
rect 2222 12180 2228 12192
rect 2280 12180 2286 12232
rect 2682 12220 2688 12232
rect 2424 12192 2688 12220
rect 2038 12112 2044 12164
rect 2096 12152 2102 12164
rect 2424 12161 2452 12192
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12220 3295 12223
rect 4154 12220 4160 12232
rect 3283 12192 4160 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 2409 12155 2467 12161
rect 2409 12152 2421 12155
rect 2096 12124 2421 12152
rect 2096 12112 2102 12124
rect 2409 12121 2421 12124
rect 2455 12121 2467 12155
rect 4724 12152 4752 12251
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 5920 12260 6009 12288
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5074 12220 5080 12232
rect 5031 12192 5080 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5684 12192 5825 12220
rect 5684 12180 5690 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 5920 12152 5948 12260
rect 5997 12257 6009 12260
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12288 6699 12291
rect 7374 12288 7380 12300
rect 6687 12260 7380 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7837 12291 7895 12297
rect 7837 12288 7849 12291
rect 7484 12260 7849 12288
rect 6822 12220 6828 12232
rect 6783 12192 6828 12220
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7484 12220 7512 12260
rect 7837 12257 7849 12260
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 9585 12291 9643 12297
rect 9585 12257 9597 12291
rect 9631 12288 9643 12291
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 9631 12260 10333 12288
rect 9631 12257 9643 12260
rect 9585 12251 9643 12257
rect 10321 12257 10333 12260
rect 10367 12288 10379 12291
rect 10962 12288 10968 12300
rect 10367 12260 10968 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 12124 12260 12541 12288
rect 12124 12248 12130 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12288 12955 12291
rect 12943 12260 13952 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13924 12232 13952 12260
rect 14642 12248 14648 12300
rect 14700 12288 14706 12300
rect 15028 12288 15056 12387
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 17954 12356 17960 12368
rect 17328 12328 17960 12356
rect 17328 12297 17356 12328
rect 17954 12316 17960 12328
rect 18012 12316 18018 12368
rect 14700 12260 14745 12288
rect 14844 12260 15056 12288
rect 17313 12291 17371 12297
rect 14700 12248 14706 12260
rect 7340 12192 7512 12220
rect 7745 12223 7803 12229
rect 7340 12180 7346 12192
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8110 12220 8116 12232
rect 7791 12192 8116 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 9306 12220 9312 12232
rect 9267 12192 9312 12220
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9824 12192 10180 12220
rect 9824 12180 9830 12192
rect 10152 12161 10180 12192
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10284 12192 10329 12220
rect 10284 12180 10290 12192
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 13044 12192 13185 12220
rect 13044 12180 13050 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 13906 12180 13912 12232
rect 13964 12180 13970 12232
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 14056 12192 14473 12220
rect 14056 12180 14062 12192
rect 14461 12189 14473 12192
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 14844 12220 14872 12260
rect 17313 12257 17325 12291
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 17586 12288 17592 12300
rect 17543 12260 17592 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 14608 12192 14872 12220
rect 15028 12192 16313 12220
rect 14608 12180 14614 12192
rect 6733 12155 6791 12161
rect 4724 12124 6684 12152
rect 2409 12115 2467 12121
rect 2774 12084 2780 12096
rect 2735 12056 2780 12084
rect 2774 12044 2780 12056
rect 2832 12044 2838 12096
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3329 12087 3387 12093
rect 2924 12056 2969 12084
rect 2924 12044 2930 12056
rect 3329 12053 3341 12087
rect 3375 12084 3387 12087
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3375 12056 3801 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4157 12087 4215 12093
rect 4157 12084 4169 12087
rect 4120 12056 4169 12084
rect 4120 12044 4126 12056
rect 4157 12053 4169 12056
rect 4203 12053 4215 12087
rect 4157 12047 4215 12053
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 4798 12084 4804 12096
rect 4295 12056 4804 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 5353 12087 5411 12093
rect 5353 12084 5365 12087
rect 5316 12056 5365 12084
rect 5316 12044 5322 12056
rect 5353 12053 5365 12056
rect 5399 12053 5411 12087
rect 5353 12047 5411 12053
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12084 5503 12087
rect 5718 12084 5724 12096
rect 5491 12056 5724 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 5905 12087 5963 12093
rect 5905 12084 5917 12087
rect 5868 12056 5917 12084
rect 5868 12044 5874 12056
rect 5905 12053 5917 12056
rect 5951 12084 5963 12087
rect 6273 12087 6331 12093
rect 6273 12084 6285 12087
rect 5951 12056 6285 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 6273 12053 6285 12056
rect 6319 12053 6331 12087
rect 6656 12084 6684 12124
rect 6733 12121 6745 12155
rect 6779 12152 6791 12155
rect 10137 12155 10195 12161
rect 6779 12124 7328 12152
rect 6779 12121 6791 12124
rect 6733 12115 6791 12121
rect 7006 12084 7012 12096
rect 6656 12056 7012 12084
rect 6273 12047 6331 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7190 12084 7196 12096
rect 7151 12056 7196 12084
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7300 12093 7328 12124
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10410 12152 10416 12164
rect 10183 12124 10416 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 12437 12155 12495 12161
rect 12437 12152 12449 12155
rect 11808 12124 12449 12152
rect 11808 12096 11836 12124
rect 12437 12121 12449 12124
rect 12483 12121 12495 12155
rect 12437 12115 12495 12121
rect 13081 12155 13139 12161
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 13127 12124 14136 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 7285 12087 7343 12093
rect 7285 12053 7297 12087
rect 7331 12053 7343 12087
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7285 12047 7343 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8536 12056 8953 12084
rect 8536 12044 8542 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 9401 12087 9459 12093
rect 9401 12084 9413 12087
rect 9272 12056 9413 12084
rect 9272 12044 9278 12056
rect 9401 12053 9413 12056
rect 9447 12053 9459 12087
rect 9766 12084 9772 12096
rect 9727 12056 9772 12084
rect 9401 12047 9459 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 11790 12084 11796 12096
rect 11751 12056 11796 12084
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12618 12084 12624 12096
rect 12391 12056 12624 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12618 12044 12624 12056
rect 12676 12084 12682 12096
rect 13354 12084 13360 12096
rect 12676 12056 13360 12084
rect 12676 12044 12682 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13538 12084 13544 12096
rect 13499 12056 13544 12084
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 13814 12084 13820 12096
rect 13775 12056 13820 12084
rect 13814 12044 13820 12056
rect 13872 12084 13878 12096
rect 13998 12084 14004 12096
rect 13872 12056 14004 12084
rect 13872 12044 13878 12056
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 14108 12093 14136 12124
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 15028 12152 15056 12192
rect 16301 12189 16313 12192
rect 16347 12220 16359 12223
rect 17678 12220 17684 12232
rect 16347 12192 17356 12220
rect 17639 12192 17684 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 14240 12124 15056 12152
rect 14240 12112 14246 12124
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 16482 12152 16488 12164
rect 16172 12124 16488 12152
rect 16172 12112 16178 12124
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 14093 12087 14151 12093
rect 14093 12053 14105 12087
rect 14139 12053 14151 12087
rect 15930 12084 15936 12096
rect 15891 12056 15936 12084
rect 14093 12047 14151 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16080 12056 16125 12084
rect 16080 12044 16086 12056
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 16577 12087 16635 12093
rect 16577 12084 16589 12087
rect 16356 12056 16589 12084
rect 16356 12044 16362 12056
rect 16577 12053 16589 12056
rect 16623 12053 16635 12087
rect 16577 12047 16635 12053
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 17126 12084 17132 12096
rect 16899 12056 17132 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 17328 12084 17356 12192
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17954 12220 17960 12232
rect 17915 12192 17960 12220
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 17770 12084 17776 12096
rect 17267 12056 17776 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2590 11880 2596 11892
rect 2551 11852 2596 11880
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 3878 11880 3884 11892
rect 3007 11852 3884 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4062 11880 4068 11892
rect 4023 11852 4068 11880
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4893 11883 4951 11889
rect 4893 11849 4905 11883
rect 4939 11880 4951 11883
rect 5074 11880 5080 11892
rect 4939 11852 5080 11880
rect 4939 11849 4951 11852
rect 4893 11843 4951 11849
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5316 11852 5457 11880
rect 5316 11840 5322 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5718 11880 5724 11892
rect 5583 11852 5724 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 6328 11852 6469 11880
rect 6328 11840 6334 11852
rect 6457 11849 6469 11852
rect 6503 11880 6515 11883
rect 7098 11880 7104 11892
rect 6503 11852 7104 11880
rect 6503 11849 6515 11852
rect 6457 11843 6515 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7285 11883 7343 11889
rect 7285 11849 7297 11883
rect 7331 11880 7343 11883
rect 7650 11880 7656 11892
rect 7331 11852 7656 11880
rect 7331 11849 7343 11852
rect 7285 11843 7343 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 8478 11880 8484 11892
rect 7800 11852 7845 11880
rect 8439 11852 8484 11880
rect 7800 11840 7806 11852
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8573 11883 8631 11889
rect 8573 11849 8585 11883
rect 8619 11880 8631 11883
rect 9766 11880 9772 11892
rect 8619 11852 9772 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10781 11883 10839 11889
rect 10781 11849 10793 11883
rect 10827 11880 10839 11883
rect 11974 11880 11980 11892
rect 10827 11852 11980 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 12360 11852 15761 11880
rect 4982 11812 4988 11824
rect 1504 11784 4988 11812
rect 1504 11756 1532 11784
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 5810 11772 5816 11824
rect 5868 11812 5874 11824
rect 9214 11812 9220 11824
rect 5868 11784 9220 11812
rect 5868 11772 5874 11784
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 9490 11812 9496 11824
rect 9324 11784 9496 11812
rect 9324 11756 9352 11784
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 9674 11772 9680 11824
rect 9732 11812 9738 11824
rect 10137 11815 10195 11821
rect 10137 11812 10149 11815
rect 9732 11784 10149 11812
rect 9732 11772 9738 11784
rect 10137 11781 10149 11784
rect 10183 11812 10195 11815
rect 10689 11815 10747 11821
rect 10689 11812 10701 11815
rect 10183 11784 10701 11812
rect 10183 11781 10195 11784
rect 10137 11775 10195 11781
rect 10689 11781 10701 11784
rect 10735 11781 10747 11815
rect 10689 11775 10747 11781
rect 11885 11815 11943 11821
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 12360 11812 12388 11852
rect 15749 11849 15761 11852
rect 15795 11849 15807 11883
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 15749 11843 15807 11849
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 11931 11784 12388 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 1486 11744 1492 11756
rect 1447 11716 1492 11744
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 1670 11704 1676 11756
rect 1728 11744 1734 11756
rect 2133 11747 2191 11753
rect 2133 11744 2145 11747
rect 1728 11716 2145 11744
rect 1728 11704 1734 11716
rect 2133 11713 2145 11716
rect 2179 11713 2191 11747
rect 3421 11747 3479 11753
rect 3421 11744 3433 11747
rect 2133 11707 2191 11713
rect 3068 11716 3433 11744
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 1118 11500 1124 11552
rect 1176 11540 1182 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 1176 11512 1593 11540
rect 1176 11500 1182 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1964 11540 1992 11639
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2096 11648 2141 11676
rect 2332 11648 2636 11676
rect 2096 11636 2102 11648
rect 2130 11568 2136 11620
rect 2188 11608 2194 11620
rect 2332 11608 2360 11648
rect 2498 11608 2504 11620
rect 2188 11580 2360 11608
rect 2459 11580 2504 11608
rect 2188 11568 2194 11580
rect 2498 11568 2504 11580
rect 2556 11568 2562 11620
rect 2608 11608 2636 11648
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3068 11685 3096 11716
rect 3421 11713 3433 11716
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11744 3939 11747
rect 4154 11744 4160 11756
rect 3927 11716 4160 11744
rect 3927 11713 3939 11716
rect 3881 11707 3939 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4356 11716 4445 11744
rect 3053 11679 3111 11685
rect 3053 11676 3065 11679
rect 2832 11648 3065 11676
rect 2832 11636 2838 11648
rect 3053 11645 3065 11648
rect 3099 11645 3111 11679
rect 3053 11639 3111 11645
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11676 3295 11679
rect 3510 11676 3516 11688
rect 3283 11648 3516 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 4356 11676 4384 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 6638 11744 6644 11756
rect 4479 11716 6644 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7156 11716 7665 11744
rect 7156 11704 7162 11716
rect 7653 11713 7665 11716
rect 7699 11744 7711 11747
rect 9306 11744 9312 11756
rect 7699 11716 9076 11744
rect 9267 11716 9312 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 4522 11676 4528 11688
rect 4172 11648 4384 11676
rect 4483 11648 4528 11676
rect 4172 11620 4200 11648
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 5353 11679 5411 11685
rect 4764 11648 4857 11676
rect 4764 11636 4770 11648
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 6086 11676 6092 11688
rect 5399 11648 6092 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6788 11648 7021 11676
rect 6788 11636 6794 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7009 11639 7067 11645
rect 7668 11648 7849 11676
rect 3697 11611 3755 11617
rect 3697 11608 3709 11611
rect 2608 11580 3709 11608
rect 3697 11577 3709 11580
rect 3743 11577 3755 11611
rect 3697 11571 3755 11577
rect 4154 11568 4160 11620
rect 4212 11568 4218 11620
rect 4246 11568 4252 11620
rect 4304 11608 4310 11620
rect 4724 11608 4752 11636
rect 6546 11608 6552 11620
rect 4304 11580 6552 11608
rect 4304 11568 4310 11580
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7098 11608 7104 11620
rect 6972 11580 7104 11608
rect 6972 11568 6978 11580
rect 7098 11568 7104 11580
rect 7156 11608 7162 11620
rect 7668 11608 7696 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 8754 11676 8760 11688
rect 8715 11648 8760 11676
rect 7837 11639 7895 11645
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 7156 11580 7696 11608
rect 7156 11568 7162 11580
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 8941 11611 8999 11617
rect 8941 11608 8953 11611
rect 7800 11580 8953 11608
rect 7800 11568 7806 11580
rect 8941 11577 8953 11580
rect 8987 11577 8999 11611
rect 9048 11608 9076 11716
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 11900 11744 11928 11775
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 14182 11812 14188 11824
rect 12492 11784 14188 11812
rect 12492 11772 12498 11784
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 14550 11772 14556 11824
rect 14608 11812 14614 11824
rect 15289 11815 15347 11821
rect 15289 11812 15301 11815
rect 14608 11784 15301 11812
rect 14608 11772 14614 11784
rect 15289 11781 15301 11784
rect 15335 11812 15347 11815
rect 15335 11784 17172 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 13446 11744 13452 11756
rect 9640 11716 10732 11744
rect 9640 11704 9646 11716
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 9272 11648 9413 11676
rect 9272 11636 9278 11648
rect 9401 11645 9413 11648
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 10134 11676 10140 11688
rect 9548 11648 9593 11676
rect 9646 11648 10140 11676
rect 9548 11636 9554 11648
rect 9646 11608 9674 11648
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 10410 11608 10416 11620
rect 9048 11580 9674 11608
rect 9784 11580 10416 11608
rect 8941 11571 8999 11577
rect 3510 11540 3516 11552
rect 1964 11512 3516 11540
rect 1581 11503 1639 11509
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 3605 11543 3663 11549
rect 3605 11509 3617 11543
rect 3651 11540 3663 11543
rect 4062 11540 4068 11552
rect 3651 11512 4068 11540
rect 3651 11509 3663 11512
rect 3605 11503 3663 11509
rect 4062 11500 4068 11512
rect 4120 11540 4126 11552
rect 5074 11540 5080 11552
rect 4120 11512 5080 11540
rect 4120 11500 4126 11512
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6181 11543 6239 11549
rect 6181 11509 6193 11543
rect 6227 11540 6239 11543
rect 6362 11540 6368 11552
rect 6227 11512 6368 11540
rect 6227 11509 6239 11512
rect 6181 11503 6239 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 6822 11540 6828 11552
rect 6735 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11540 6886 11552
rect 7926 11540 7932 11552
rect 6880 11512 7932 11540
rect 6880 11500 6886 11512
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8386 11540 8392 11552
rect 8159 11512 8392 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9784 11549 9812 11580
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 10704 11608 10732 11716
rect 11072 11716 11928 11744
rect 13407 11716 13452 11744
rect 10962 11676 10968 11688
rect 10923 11648 10968 11676
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11072 11608 11100 11716
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13630 11744 13636 11756
rect 13556 11716 13636 11744
rect 11974 11676 11980 11688
rect 11935 11648 11980 11676
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12124 11648 12217 11676
rect 12124 11636 12130 11648
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 13556 11685 13584 11716
rect 13630 11704 13636 11716
rect 13688 11744 13694 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13688 11716 13921 11744
rect 13688 11704 13694 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 14918 11704 14924 11756
rect 14976 11744 14982 11756
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 14976 11716 15209 11744
rect 14976 11704 14982 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 12768 11648 13553 11676
rect 12768 11636 12774 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13722 11676 13728 11688
rect 13683 11648 13728 11676
rect 13541 11639 13599 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11645 15163 11679
rect 15212 11676 15240 11707
rect 15948 11676 15976 11707
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16908 11716 17049 11744
rect 16908 11704 16914 11716
rect 17037 11713 17049 11716
rect 17083 11713 17095 11747
rect 17144 11744 17172 11784
rect 17218 11772 17224 11824
rect 17276 11812 17282 11824
rect 17276 11784 18460 11812
rect 17276 11772 17282 11784
rect 18432 11756 18460 11784
rect 17494 11744 17500 11756
rect 17144 11716 17500 11744
rect 17037 11707 17095 11713
rect 17494 11704 17500 11716
rect 17552 11744 17558 11756
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 17552 11716 17601 11744
rect 17552 11704 17558 11716
rect 17589 11713 17601 11716
rect 17635 11713 17647 11747
rect 18046 11744 18052 11756
rect 18007 11716 18052 11744
rect 17589 11707 17647 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 15212 11648 15976 11676
rect 15105 11639 15163 11645
rect 10704 11580 11100 11608
rect 11238 11568 11244 11620
rect 11296 11608 11302 11620
rect 12084 11608 12112 11636
rect 14550 11608 14556 11620
rect 11296 11580 12112 11608
rect 14511 11580 14556 11608
rect 11296 11568 11302 11580
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 15120 11608 15148 11639
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 16264 11648 16405 11676
rect 16264 11636 16270 11648
rect 16393 11645 16405 11648
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 17126 11676 17132 11688
rect 16540 11648 17132 11676
rect 16540 11636 16546 11648
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 15838 11608 15844 11620
rect 15120 11580 15844 11608
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 17236 11608 17264 11639
rect 15948 11580 17264 11608
rect 17773 11611 17831 11617
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9364 11512 9781 11540
rect 9364 11500 9370 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 9769 11503 9827 11509
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9916 11512 10333 11540
rect 9916 11500 9922 11512
rect 10321 11509 10333 11512
rect 10367 11509 10379 11543
rect 10321 11503 10379 11509
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 10560 11512 11529 11540
rect 10560 11500 10566 11512
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 11517 11503 11575 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14734 11540 14740 11552
rect 14424 11512 14740 11540
rect 14424 11500 14430 11512
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 15657 11543 15715 11549
rect 15657 11540 15669 11543
rect 15528 11512 15669 11540
rect 15528 11500 15534 11512
rect 15657 11509 15669 11512
rect 15703 11509 15715 11543
rect 15657 11503 15715 11509
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 15948 11540 15976 11580
rect 17773 11577 17785 11611
rect 17819 11608 17831 11611
rect 18690 11608 18696 11620
rect 17819 11580 18696 11608
rect 17819 11577 17831 11580
rect 17773 11571 17831 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 16114 11540 16120 11552
rect 15804 11512 15976 11540
rect 16075 11512 16120 11540
rect 15804 11500 15810 11512
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11540 16359 11543
rect 16390 11540 16396 11552
rect 16347 11512 16396 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16669 11543 16727 11549
rect 16669 11509 16681 11543
rect 16715 11540 16727 11543
rect 16942 11540 16948 11552
rect 16715 11512 16948 11540
rect 16715 11509 16727 11512
rect 16669 11503 16727 11509
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 17957 11543 18015 11549
rect 17957 11540 17969 11543
rect 17920 11512 17969 11540
rect 17920 11500 17926 11512
rect 17957 11509 17969 11512
rect 18003 11509 18015 11543
rect 17957 11503 18015 11509
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 18288 11512 18337 11540
rect 18288 11500 18294 11512
rect 18325 11509 18337 11512
rect 18371 11509 18383 11543
rect 18325 11503 18383 11509
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 1820 11308 3525 11336
rect 1820 11296 1826 11308
rect 3513 11305 3525 11308
rect 3559 11336 3571 11339
rect 3786 11336 3792 11348
rect 3559 11308 3792 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4525 11339 4583 11345
rect 3896 11308 4476 11336
rect 1854 11228 1860 11280
rect 1912 11268 1918 11280
rect 2317 11271 2375 11277
rect 2317 11268 2329 11271
rect 1912 11240 2329 11268
rect 1912 11228 1918 11240
rect 2317 11237 2329 11240
rect 2363 11237 2375 11271
rect 2317 11231 2375 11237
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 3896 11268 3924 11308
rect 4154 11268 4160 11280
rect 3467 11240 3924 11268
rect 4080 11240 4160 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 2406 11160 2412 11212
rect 2464 11200 2470 11212
rect 4080 11209 4108 11240
rect 4154 11228 4160 11240
rect 4212 11228 4218 11280
rect 4448 11268 4476 11308
rect 4525 11305 4537 11339
rect 4571 11336 4583 11339
rect 4798 11336 4804 11348
rect 4571 11308 4804 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 7558 11336 7564 11348
rect 6696 11308 7564 11336
rect 6696 11296 6702 11308
rect 7558 11296 7564 11308
rect 7616 11336 7622 11348
rect 8570 11336 8576 11348
rect 7616 11308 8576 11336
rect 7616 11296 7622 11308
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 11054 11336 11060 11348
rect 8803 11308 11060 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 15010 11336 15016 11348
rect 14971 11308 15016 11336
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15378 11296 15384 11348
rect 15436 11336 15442 11348
rect 16390 11336 16396 11348
rect 15436 11308 16396 11336
rect 15436 11296 15442 11308
rect 16390 11296 16396 11308
rect 16448 11336 16454 11348
rect 16850 11336 16856 11348
rect 16448 11308 16712 11336
rect 16811 11308 16856 11336
rect 16448 11296 16454 11308
rect 4448 11240 4752 11268
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 2464 11172 2789 11200
rect 2464 11160 2470 11172
rect 2777 11169 2789 11172
rect 2823 11169 2835 11203
rect 2777 11163 2835 11169
rect 3881 11203 3939 11209
rect 3881 11169 3893 11203
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11169 4123 11203
rect 4246 11200 4252 11212
rect 4065 11163 4123 11169
rect 4172 11172 4252 11200
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11101 2007 11135
rect 2222 11132 2228 11144
rect 2183 11104 2228 11132
rect 1949 11095 2007 11101
rect 1964 10996 1992 11095
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3896 11132 3924 11163
rect 4172 11132 4200 11172
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 3896 11104 4200 11132
rect 4724 11132 4752 11240
rect 4890 11228 4896 11280
rect 4948 11268 4954 11280
rect 5537 11271 5595 11277
rect 5537 11268 5549 11271
rect 4948 11240 5549 11268
rect 4948 11228 4954 11240
rect 5537 11237 5549 11240
rect 5583 11237 5595 11271
rect 6365 11271 6423 11277
rect 5537 11231 5595 11237
rect 5828 11240 6224 11268
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 5828 11200 5856 11240
rect 5994 11200 6000 11212
rect 4847 11172 5856 11200
rect 5955 11172 6000 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6196 11209 6224 11240
rect 6365 11237 6377 11271
rect 6411 11237 6423 11271
rect 7466 11268 7472 11280
rect 6365 11231 6423 11237
rect 6932 11240 7472 11268
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11200 6239 11203
rect 6270 11200 6276 11212
rect 6227 11172 6276 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4724 11104 4997 11132
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 6380 11132 6408 11231
rect 6932 11209 6960 11240
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 9309 11271 9367 11277
rect 9309 11268 9321 11271
rect 8496 11240 9321 11268
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 5951 11104 6408 11132
rect 6472 11172 6929 11200
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2740 11036 2973 11064
rect 2740 11024 2746 11036
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 2961 11027 3019 11033
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4028 11036 4905 11064
rect 4028 11024 4034 11036
rect 4893 11033 4905 11036
rect 4939 11033 4951 11067
rect 6472 11064 6500 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 7650 11200 7656 11212
rect 7064 11172 7656 11200
rect 7064 11160 7070 11172
rect 7650 11160 7656 11172
rect 7708 11200 7714 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7708 11172 7757 11200
rect 7708 11160 7714 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11200 8355 11203
rect 8496 11200 8524 11240
rect 9309 11237 9321 11240
rect 9355 11237 9367 11271
rect 10410 11268 10416 11280
rect 9309 11231 9367 11237
rect 9646 11240 10416 11268
rect 8343 11172 8524 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7558 11132 7564 11144
rect 6880 11104 6925 11132
rect 7519 11104 7564 11132
rect 6880 11092 6886 11104
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 6546 11064 6552 11076
rect 4893 11027 4951 11033
rect 5000 11036 6552 11064
rect 5000 11008 5028 11036
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 7282 11064 7288 11076
rect 6972 11036 7288 11064
rect 6972 11024 6978 11036
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7653 11067 7711 11073
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 8220 11064 8248 11163
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 9646 11200 9674 11240
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 10965 11271 11023 11277
rect 10965 11268 10977 11271
rect 10520 11240 10977 11268
rect 8628 11172 9674 11200
rect 9861 11203 9919 11209
rect 8628 11160 8634 11172
rect 9861 11169 9873 11203
rect 9907 11169 9919 11203
rect 10520 11200 10548 11240
rect 10965 11237 10977 11240
rect 11011 11237 11023 11271
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 10965 11231 11023 11237
rect 13004 11240 14105 11268
rect 9861 11163 9919 11169
rect 10336 11172 10548 11200
rect 10781 11203 10839 11209
rect 8386 11132 8392 11144
rect 8347 11104 8392 11132
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9582 11132 9588 11144
rect 8680 11104 9588 11132
rect 8478 11064 8484 11076
rect 7699 11036 8187 11064
rect 8220 11036 8484 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 3142 10996 3148 11008
rect 1964 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 4157 10999 4215 11005
rect 4157 10965 4169 10999
rect 4203 10996 4215 10999
rect 4246 10996 4252 11008
rect 4203 10968 4252 10996
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 4982 10956 4988 11008
rect 5040 10956 5046 11008
rect 5258 10956 5264 11008
rect 5316 10996 5322 11008
rect 5353 10999 5411 11005
rect 5353 10996 5365 10999
rect 5316 10968 5365 10996
rect 5316 10956 5322 10968
rect 5353 10965 5365 10968
rect 5399 10965 5411 10999
rect 7190 10996 7196 11008
rect 7151 10968 7196 10996
rect 5353 10959 5411 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 8159 10996 8187 11036
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 8680 10996 8708 11104
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9732 11104 9777 11132
rect 9732 11092 9738 11104
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 9876 11064 9904 11163
rect 8812 11036 9904 11064
rect 10336 11064 10364 11172
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 10502 11132 10508 11144
rect 10463 11104 10508 11132
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10612 11064 10640 11095
rect 10336 11036 10640 11064
rect 8812 11024 8818 11036
rect 8938 10996 8944 11008
rect 8159 10968 8708 10996
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9214 10996 9220 11008
rect 9175 10968 9220 10996
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9769 10999 9827 11005
rect 9769 10965 9781 10999
rect 9815 10996 9827 10999
rect 10137 10999 10195 11005
rect 10137 10996 10149 10999
rect 9815 10968 10149 10996
rect 9815 10965 9827 10968
rect 9769 10959 9827 10965
rect 10137 10965 10149 10968
rect 10183 10965 10195 10999
rect 10137 10959 10195 10965
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 10796 10996 10824 11163
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 13004 11209 13032 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 16577 11271 16635 11277
rect 16577 11268 16589 11271
rect 14976 11240 16589 11268
rect 14976 11228 14982 11240
rect 16577 11237 16589 11240
rect 16623 11237 16635 11271
rect 16684 11268 16712 11308
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 18966 11268 18972 11280
rect 16684 11240 18972 11268
rect 16577 11231 16635 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11296 11172 11529 11200
rect 11296 11160 11302 11172
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 11333 11067 11391 11073
rect 11333 11033 11345 11067
rect 11379 11064 11391 11067
rect 11514 11064 11520 11076
rect 11379 11036 11520 11064
rect 11379 11033 11391 11036
rect 11333 11027 11391 11033
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 12912 11064 12940 11163
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 13504 11172 13553 11200
rect 13504 11160 13510 11172
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 13541 11163 13599 11169
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 13780 11172 14657 11200
rect 13780 11160 13786 11172
rect 14645 11169 14657 11172
rect 14691 11200 14703 11203
rect 15562 11200 15568 11212
rect 14691 11172 15568 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15746 11200 15752 11212
rect 15707 11172 15752 11200
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 15930 11160 15936 11212
rect 15988 11200 15994 11212
rect 15988 11172 16896 11200
rect 15988 11160 15994 11172
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 14366 11132 14372 11144
rect 13228 11104 14372 11132
rect 13228 11092 13234 11104
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 14424 11104 14565 11132
rect 14424 11092 14430 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 15470 11132 15476 11144
rect 15431 11104 15476 11132
rect 14553 11095 14611 11101
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 16206 11132 16212 11144
rect 16167 11104 16212 11132
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 16298 11092 16304 11144
rect 16356 11132 16362 11144
rect 16356 11104 16401 11132
rect 16356 11092 16362 11104
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 16761 11135 16819 11141
rect 16761 11132 16773 11135
rect 16632 11104 16773 11132
rect 16632 11092 16638 11104
rect 16761 11101 16773 11104
rect 16807 11101 16819 11135
rect 16868 11132 16896 11172
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 17313 11203 17371 11209
rect 17313 11200 17325 11203
rect 17184 11172 17325 11200
rect 17184 11160 17190 11172
rect 17313 11169 17325 11172
rect 17359 11169 17371 11203
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 17313 11163 17371 11169
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 17678 11132 17684 11144
rect 16868 11104 17684 11132
rect 16761 11095 16819 11101
rect 13722 11064 13728 11076
rect 12912 11036 13728 11064
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 13872 11036 14473 11064
rect 13872 11024 13878 11036
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 15565 11067 15623 11073
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 16666 11064 16672 11076
rect 15611 11036 16672 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 16776 11064 16804 11095
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17954 11132 17960 11144
rect 17915 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 17402 11064 17408 11076
rect 16776 11036 17408 11064
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 10962 10996 10968 11008
rect 10652 10968 10968 10996
rect 10652 10956 10658 10968
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 11425 10999 11483 11005
rect 11425 10965 11437 10999
rect 11471 10996 11483 10999
rect 11790 10996 11796 11008
rect 11471 10968 11796 10996
rect 11471 10965 11483 10968
rect 11425 10959 11483 10965
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 13446 10996 13452 11008
rect 13407 10968 13452 10996
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 15102 10996 15108 11008
rect 15063 10968 15108 10996
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 15930 10956 15936 11008
rect 15988 10996 15994 11008
rect 16025 10999 16083 11005
rect 16025 10996 16037 10999
rect 15988 10968 16037 10996
rect 15988 10956 15994 10968
rect 16025 10965 16037 10968
rect 16071 10965 16083 10999
rect 16025 10959 16083 10965
rect 16485 10999 16543 11005
rect 16485 10965 16497 10999
rect 16531 10996 16543 10999
rect 17034 10996 17040 11008
rect 16531 10968 17040 10996
rect 16531 10965 16543 10968
rect 16485 10959 16543 10965
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 17218 10996 17224 11008
rect 17179 10968 17224 10996
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 1946 10752 1952 10804
rect 2004 10792 2010 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 2004 10764 2053 10792
rect 2004 10752 2010 10764
rect 2041 10761 2053 10764
rect 2087 10792 2099 10795
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2087 10764 2513 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2501 10755 2559 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3050 10792 3056 10804
rect 2963 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10792 3114 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3108 10764 3617 10792
rect 3108 10752 3114 10764
rect 3605 10761 3617 10764
rect 3651 10792 3663 10795
rect 3651 10764 3924 10792
rect 3651 10761 3663 10764
rect 3605 10755 3663 10761
rect 2222 10684 2228 10736
rect 2280 10724 2286 10736
rect 3896 10733 3924 10764
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 4028 10764 4077 10792
rect 4028 10752 4034 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4522 10792 4528 10804
rect 4295 10764 4528 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5810 10792 5816 10804
rect 5040 10764 5816 10792
rect 5040 10752 5046 10764
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6362 10792 6368 10804
rect 5951 10764 6368 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 8846 10792 8852 10804
rect 6656 10764 8852 10792
rect 3697 10727 3755 10733
rect 3697 10724 3709 10727
rect 2280 10696 3709 10724
rect 2280 10684 2286 10696
rect 3697 10693 3709 10696
rect 3743 10693 3755 10727
rect 3697 10687 3755 10693
rect 3881 10727 3939 10733
rect 3881 10693 3893 10727
rect 3927 10724 3939 10727
rect 4617 10727 4675 10733
rect 4617 10724 4629 10727
rect 3927 10696 4629 10724
rect 3927 10693 3939 10696
rect 3881 10687 3939 10693
rect 4617 10693 4629 10696
rect 4663 10724 4675 10727
rect 4663 10696 5856 10724
rect 4663 10693 4675 10696
rect 4617 10687 4675 10693
rect 5828 10668 5856 10696
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10625 1639 10659
rect 2314 10656 2320 10668
rect 1581 10619 1639 10625
rect 1780 10628 2320 10656
rect 1596 10520 1624 10619
rect 1780 10597 1808 10628
rect 2314 10616 2320 10628
rect 2372 10656 2378 10668
rect 2682 10656 2688 10668
rect 2372 10628 2688 10656
rect 2372 10616 2378 10628
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 4982 10656 4988 10668
rect 3200 10628 4988 10656
rect 3200 10616 3206 10628
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1765 10551 1823 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3510 10588 3516 10600
rect 3375 10560 3516 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 4724 10597 4752 10628
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 5224 10628 5273 10656
rect 5224 10616 5230 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6236 10628 6561 10656
rect 6236 10616 6242 10628
rect 6549 10625 6561 10628
rect 6595 10656 6607 10659
rect 6656 10656 6684 10764
rect 8846 10752 8852 10764
rect 8904 10752 8910 10804
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 12618 10792 12624 10804
rect 10284 10764 12624 10792
rect 10284 10752 10290 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 12894 10792 12900 10804
rect 12855 10764 12900 10792
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 13446 10792 13452 10804
rect 13311 10764 13452 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 15102 10792 15108 10804
rect 14507 10764 15108 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 15252 10764 15297 10792
rect 15488 10764 15761 10792
rect 15252 10752 15258 10764
rect 6917 10727 6975 10733
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 11974 10724 11980 10736
rect 6963 10696 11980 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 13630 10724 13636 10736
rect 13280 10696 13636 10724
rect 6595 10628 6684 10656
rect 6733 10659 6791 10665
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6779 10628 7389 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 8251 10628 9597 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 4709 10591 4767 10597
rect 4709 10557 4721 10591
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 3050 10520 3056 10532
rect 1596 10492 3056 10520
rect 3050 10480 3056 10492
rect 3108 10480 3114 10532
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 4816 10520 4844 10551
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5626 10588 5632 10600
rect 5132 10560 5632 10588
rect 5132 10548 5138 10560
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6454 10588 6460 10600
rect 6135 10560 6460 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 6748 10520 6776 10619
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 9824 10628 10517 10656
rect 9824 10616 9830 10628
rect 10505 10625 10517 10628
rect 10551 10656 10563 10659
rect 10962 10656 10968 10668
rect 10551 10628 10968 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11330 10656 11336 10668
rect 11291 10628 11336 10656
rect 11330 10616 11336 10628
rect 11388 10656 11394 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11388 10628 11897 10656
rect 11388 10616 11394 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 13280 10656 13308 10696
rect 13630 10684 13636 10696
rect 13688 10724 13694 10736
rect 13814 10724 13820 10736
rect 13688 10696 13820 10724
rect 13688 10684 13694 10696
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14369 10727 14427 10733
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 14734 10724 14740 10736
rect 14415 10696 14740 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 11931 10628 13308 10656
rect 13357 10659 13415 10665
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 14182 10656 14188 10668
rect 13403 10628 14188 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 15488 10656 15516 10764
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 16172 10764 16221 10792
rect 16172 10752 16178 10764
rect 16209 10761 16221 10764
rect 16255 10761 16267 10795
rect 16666 10792 16672 10804
rect 16627 10764 16672 10792
rect 16209 10755 16267 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 16776 10764 17172 10792
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 16776 10724 16804 10764
rect 15896 10696 16804 10724
rect 15896 10684 15902 10696
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15335 10628 15516 10656
rect 15580 10628 16129 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7006 10588 7012 10600
rect 6880 10560 7012 10588
rect 6880 10548 6886 10560
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10557 7527 10591
rect 7650 10588 7656 10600
rect 7611 10560 7656 10588
rect 7469 10551 7527 10557
rect 4580 10492 4844 10520
rect 5092 10492 6776 10520
rect 7484 10520 7512 10551
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10557 8355 10591
rect 8297 10551 8355 10557
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8570 10588 8576 10600
rect 8527 10560 8576 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8018 10520 8024 10532
rect 7484 10492 8024 10520
rect 4580 10480 4586 10492
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 5092 10461 5120 10492
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 5077 10455 5135 10461
rect 5077 10452 5089 10455
rect 4396 10424 5089 10452
rect 4396 10412 4402 10424
rect 5077 10421 5089 10424
rect 5123 10421 5135 10455
rect 5442 10452 5448 10464
rect 5403 10424 5448 10452
rect 5077 10415 5135 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6052 10424 6377 10452
rect 6052 10412 6058 10424
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 7006 10452 7012 10464
rect 6967 10424 7012 10452
rect 6365 10415 6423 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7524 10424 7849 10452
rect 7524 10412 7530 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 7837 10415 7895 10421
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8312 10452 8340 10551
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 8941 10591 8999 10597
rect 8720 10560 8765 10588
rect 8720 10548 8726 10560
rect 8941 10557 8953 10591
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 8956 10520 8984 10551
rect 10410 10548 10416 10600
rect 10468 10588 10474 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10468 10560 10609 10588
rect 10468 10548 10474 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 11606 10588 11612 10600
rect 10827 10560 11612 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10588 11851 10591
rect 12434 10588 12440 10600
rect 11839 10560 12440 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 11716 10520 11744 10551
rect 12434 10548 12440 10560
rect 12492 10588 12498 10600
rect 13446 10588 13452 10600
rect 12492 10560 12585 10588
rect 13407 10560 13452 10588
rect 12492 10548 12498 10560
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 13872 10560 14565 10588
rect 13872 10548 13878 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14642 10548 14648 10600
rect 14700 10588 14706 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 14700 10560 15393 10588
rect 14700 10548 14706 10560
rect 15381 10557 15393 10560
rect 15427 10588 15439 10591
rect 15470 10588 15476 10600
rect 15427 10560 15476 10588
rect 15427 10557 15439 10560
rect 15381 10551 15439 10557
rect 15470 10548 15476 10560
rect 15528 10548 15534 10600
rect 12802 10520 12808 10532
rect 8956 10492 11376 10520
rect 11716 10492 12808 10520
rect 8938 10452 8944 10464
rect 8260 10424 8944 10452
rect 8260 10412 8266 10424
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 10137 10455 10195 10461
rect 10137 10421 10149 10455
rect 10183 10452 10195 10455
rect 10226 10452 10232 10464
rect 10183 10424 10232 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10962 10452 10968 10464
rect 10923 10424 10968 10452
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11348 10452 11376 10492
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 13909 10523 13967 10529
rect 13909 10520 13921 10523
rect 13228 10492 13921 10520
rect 13228 10480 13234 10492
rect 13909 10489 13921 10492
rect 13955 10520 13967 10523
rect 15580 10520 15608 10628
rect 16117 10625 16129 10628
rect 16163 10656 16175 10659
rect 16758 10656 16764 10668
rect 16163 10628 16764 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16960 10628 17049 10656
rect 16960 10600 16988 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17144 10656 17172 10764
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17276 10764 17509 10792
rect 17276 10752 17282 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 18046 10792 18052 10804
rect 17497 10755 17555 10761
rect 17972 10764 18052 10792
rect 17144 10628 17264 10656
rect 17037 10619 17095 10625
rect 16301 10591 16359 10597
rect 16301 10588 16313 10591
rect 13955 10492 15608 10520
rect 15672 10560 16313 10588
rect 13955 10489 13967 10492
rect 13909 10483 13967 10489
rect 11790 10452 11796 10464
rect 11348 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 12032 10424 12265 10452
rect 12032 10412 12038 10424
rect 12253 10421 12265 10424
rect 12299 10421 12311 10455
rect 12618 10452 12624 10464
rect 12579 10424 12624 10452
rect 12253 10415 12311 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14516 10424 14841 10452
rect 14516 10412 14522 10424
rect 14829 10421 14841 10424
rect 14875 10421 14887 10455
rect 14829 10415 14887 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 15672 10452 15700 10560
rect 16301 10557 16313 10560
rect 16347 10557 16359 10591
rect 16301 10551 16359 10557
rect 16942 10548 16948 10600
rect 17000 10548 17006 10600
rect 17126 10588 17132 10600
rect 17087 10560 17132 10588
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17236 10588 17264 10628
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 17236 10560 17325 10588
rect 17313 10557 17325 10560
rect 17359 10588 17371 10591
rect 17494 10588 17500 10600
rect 17359 10560 17500 10588
rect 17359 10557 17371 10560
rect 17313 10551 17371 10557
rect 17494 10548 17500 10560
rect 17552 10548 17558 10600
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 17972 10588 18000 10764
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18138 10656 18144 10668
rect 18095 10628 18144 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 18233 10591 18291 10597
rect 18233 10588 18245 10591
rect 17920 10560 18245 10588
rect 17920 10548 17926 10560
rect 18233 10557 18245 10560
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 18432 10532 18460 10619
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 18414 10520 18420 10532
rect 16080 10492 18420 10520
rect 16080 10480 16086 10492
rect 18414 10480 18420 10492
rect 18472 10480 18478 10532
rect 15252 10424 15700 10452
rect 15252 10412 15258 10424
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 17034 10452 17040 10464
rect 15804 10424 17040 10452
rect 15804 10412 15810 10424
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17865 10455 17923 10461
rect 17865 10452 17877 10455
rect 17276 10424 17877 10452
rect 17276 10412 17282 10424
rect 17865 10421 17877 10424
rect 17911 10421 17923 10455
rect 17865 10415 17923 10421
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 2556 10220 2605 10248
rect 2556 10208 2562 10220
rect 2593 10217 2605 10220
rect 2639 10217 2651 10251
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 2593 10211 2651 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 3881 10251 3939 10257
rect 3881 10217 3893 10251
rect 3927 10248 3939 10251
rect 4246 10248 4252 10260
rect 3927 10220 4252 10248
rect 3927 10217 3939 10220
rect 3881 10211 3939 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4816 10220 5580 10248
rect 2409 10183 2467 10189
rect 2409 10149 2421 10183
rect 2455 10180 2467 10183
rect 4614 10180 4620 10192
rect 2455 10152 4620 10180
rect 2455 10149 2467 10152
rect 2409 10143 2467 10149
rect 2424 10112 2452 10143
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 4709 10183 4767 10189
rect 4709 10149 4721 10183
rect 4755 10149 4767 10183
rect 4709 10143 4767 10149
rect 1872 10084 2452 10112
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 1872 10053 1900 10084
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 2648 10084 3525 10112
rect 2648 10072 2654 10084
rect 3513 10081 3525 10084
rect 3559 10081 3571 10115
rect 4338 10112 4344 10124
rect 4299 10084 4344 10112
rect 3513 10075 3571 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 2498 10044 2504 10056
rect 2087 10016 2504 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 2777 10047 2835 10053
rect 2777 10044 2789 10047
rect 2740 10016 2789 10044
rect 2740 10004 2746 10016
rect 2777 10013 2789 10016
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 4724 10044 4752 10143
rect 3844 10016 4752 10044
rect 3844 10004 3850 10016
rect 1504 9976 1532 10004
rect 2222 9976 2228 9988
rect 1504 9948 2084 9976
rect 2183 9948 2228 9976
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2056 9908 2084 9948
rect 2222 9936 2228 9948
rect 2280 9976 2286 9988
rect 3329 9979 3387 9985
rect 3329 9976 3341 9979
rect 2280 9948 3341 9976
rect 2280 9936 2286 9948
rect 3329 9945 3341 9948
rect 3375 9945 3387 9979
rect 4246 9976 4252 9988
rect 4207 9948 4252 9976
rect 3329 9939 3387 9945
rect 4246 9936 4252 9948
rect 4304 9976 4310 9988
rect 4816 9976 4844 10220
rect 5350 10180 5356 10192
rect 5184 10152 5356 10180
rect 5184 10121 5212 10152
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5258 10072 5264 10124
rect 5316 10112 5322 10124
rect 5316 10084 5361 10112
rect 5316 10072 5322 10084
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5552 10044 5580 10220
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 8018 10248 8024 10260
rect 6420 10220 7788 10248
rect 7979 10220 8024 10248
rect 6420 10208 6426 10220
rect 7006 10180 7012 10192
rect 6840 10152 7012 10180
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5684 10084 6009 10112
rect 5684 10072 5690 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6638 10112 6644 10124
rect 6227 10084 6644 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 5132 10016 5177 10044
rect 5552 10016 5856 10044
rect 5132 10004 5138 10016
rect 5828 9988 5856 10016
rect 4304 9948 4844 9976
rect 5184 9948 5580 9976
rect 4304 9936 4310 9948
rect 2590 9908 2596 9920
rect 2056 9880 2596 9908
rect 2590 9868 2596 9880
rect 2648 9868 2654 9920
rect 3142 9908 3148 9920
rect 3103 9880 3148 9908
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 4338 9908 4344 9920
rect 3936 9880 4344 9908
rect 3936 9868 3942 9880
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 5184 9908 5212 9948
rect 5552 9917 5580 9948
rect 5810 9936 5816 9988
rect 5868 9936 5874 9988
rect 6012 9976 6040 10075
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6840 10121 6868 10152
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10081 6883 10115
rect 6825 10075 6883 10081
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10081 6975 10115
rect 7282 10112 7288 10124
rect 7243 10084 7288 10112
rect 6917 10075 6975 10081
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6932 10044 6960 10075
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7760 10112 7788 10220
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 11020 10220 18337 10248
rect 11020 10208 11026 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 7834 10140 7840 10192
rect 7892 10180 7898 10192
rect 8202 10180 8208 10192
rect 7892 10152 8208 10180
rect 7892 10140 7898 10152
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 9306 10180 9312 10192
rect 8312 10152 9312 10180
rect 8312 10112 8340 10152
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 11514 10180 11520 10192
rect 9692 10152 11520 10180
rect 7392 10084 7696 10112
rect 7760 10084 8340 10112
rect 6144 10016 6960 10044
rect 6144 10004 6150 10016
rect 7392 9976 7420 10084
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7524 10016 7573 10044
rect 7524 10004 7530 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7668 10044 7696 10084
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8573 10115 8631 10121
rect 8573 10112 8585 10115
rect 8444 10084 8585 10112
rect 8444 10072 8450 10084
rect 8573 10081 8585 10084
rect 8619 10081 8631 10115
rect 8938 10112 8944 10124
rect 8851 10084 8944 10112
rect 8573 10075 8631 10081
rect 8938 10072 8944 10084
rect 8996 10112 9002 10124
rect 9582 10112 9588 10124
rect 8996 10084 9588 10112
rect 8996 10072 9002 10084
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 7668 10016 8493 10044
rect 7561 10007 7619 10013
rect 8481 10013 8493 10016
rect 8527 10044 8539 10047
rect 8662 10044 8668 10056
rect 8527 10016 8668 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 8202 9976 8208 9988
rect 6012 9948 7420 9976
rect 7484 9948 8208 9976
rect 4856 9880 5212 9908
rect 5537 9911 5595 9917
rect 4856 9868 4862 9880
rect 5537 9877 5549 9911
rect 5583 9877 5595 9911
rect 5537 9871 5595 9877
rect 5905 9911 5963 9917
rect 5905 9877 5917 9911
rect 5951 9908 5963 9911
rect 6178 9908 6184 9920
rect 5951 9880 6184 9908
rect 5951 9877 5963 9880
rect 5905 9871 5963 9877
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6362 9908 6368 9920
rect 6323 9880 6368 9908
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 6733 9911 6791 9917
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 7190 9908 7196 9920
rect 6779 9880 7196 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7484 9917 7512 9948
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 9232 9976 9260 10007
rect 8352 9948 9260 9976
rect 8352 9936 8358 9948
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9877 7527 9911
rect 7926 9908 7932 9920
rect 7887 9880 7932 9908
rect 7469 9871 7527 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 8846 9908 8852 9920
rect 8435 9880 8852 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8846 9868 8852 9880
rect 8904 9908 8910 9920
rect 9692 9908 9720 10152
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 11940 10152 12434 10180
rect 11940 10140 11946 10152
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 10962 10112 10968 10124
rect 10744 10084 10968 10112
rect 10744 10072 10750 10084
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 12066 10112 12072 10124
rect 11195 10084 12072 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11882 10044 11888 10056
rect 11655 10016 11888 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 12406 10044 12434 10152
rect 12526 10140 12532 10192
rect 12584 10180 12590 10192
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 12584 10152 13093 10180
rect 12584 10140 12590 10152
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 15746 10180 15752 10192
rect 13081 10143 13139 10149
rect 13832 10152 15752 10180
rect 12802 10112 12808 10124
rect 12763 10084 12808 10112
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13044 10084 13645 10112
rect 13044 10072 13050 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 13354 10044 13360 10056
rect 12406 10016 13360 10044
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 13538 10044 13544 10056
rect 13495 10016 13544 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 12618 9976 12624 9988
rect 10919 9948 12296 9976
rect 12531 9948 12624 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 10502 9908 10508 9920
rect 8904 9880 9720 9908
rect 10463 9880 10508 9908
rect 8904 9868 8910 9880
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10965 9911 11023 9917
rect 10965 9877 10977 9911
rect 11011 9908 11023 9911
rect 11238 9908 11244 9920
rect 11011 9880 11244 9908
rect 11011 9877 11023 9880
rect 10965 9871 11023 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 12268 9917 12296 9948
rect 12618 9936 12624 9948
rect 12676 9976 12682 9988
rect 13832 9976 13860 10152
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 17586 10180 17592 10192
rect 16132 10152 16344 10180
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 13964 10084 14749 10112
rect 13964 10072 13970 10084
rect 14737 10081 14749 10084
rect 14783 10112 14795 10115
rect 15102 10112 15108 10124
rect 14783 10084 15108 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 16132 10112 16160 10152
rect 16316 10121 16344 10152
rect 17420 10152 17592 10180
rect 15620 10084 16160 10112
rect 16301 10115 16359 10121
rect 15620 10072 15626 10084
rect 16301 10081 16313 10115
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 17221 10115 17279 10121
rect 17221 10081 17233 10115
rect 17267 10112 17279 10115
rect 17420 10112 17448 10152
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 17773 10183 17831 10189
rect 17773 10149 17785 10183
rect 17819 10180 17831 10183
rect 18138 10180 18144 10192
rect 17819 10152 18144 10180
rect 17819 10149 17831 10152
rect 17773 10143 17831 10149
rect 18138 10140 18144 10152
rect 18196 10140 18202 10192
rect 17862 10112 17868 10124
rect 17267 10084 17448 10112
rect 17696 10084 17868 10112
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 14458 10044 14464 10056
rect 14419 10016 14464 10044
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 16209 10047 16267 10053
rect 15436 10016 15976 10044
rect 15436 10004 15442 10016
rect 12676 9948 13860 9976
rect 12676 9936 12682 9948
rect 12253 9911 12311 9917
rect 12253 9877 12265 9911
rect 12299 9877 12311 9911
rect 12253 9871 12311 9877
rect 12713 9911 12771 9917
rect 12713 9877 12725 9911
rect 12759 9908 12771 9911
rect 13078 9908 13084 9920
rect 12759 9880 13084 9908
rect 12759 9877 12771 9880
rect 12713 9871 12771 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13541 9911 13599 9917
rect 13541 9877 13553 9911
rect 13587 9908 13599 9911
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13587 9880 14105 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14599 9880 14933 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 14921 9871 14979 9877
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 15068 9880 15301 9908
rect 15068 9868 15074 9880
rect 15289 9877 15301 9880
rect 15335 9877 15347 9911
rect 15289 9871 15347 9877
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 15746 9908 15752 9920
rect 15436 9880 15481 9908
rect 15707 9880 15752 9908
rect 15436 9868 15442 9880
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 15948 9908 15976 10016
rect 16209 10013 16221 10047
rect 16255 10020 16267 10047
rect 16255 10013 16436 10020
rect 16209 10007 16436 10013
rect 16224 9992 16436 10007
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17402 10044 17408 10056
rect 17092 10016 17408 10044
rect 17092 10004 17098 10016
rect 17402 10004 17408 10016
rect 17460 10044 17466 10056
rect 17589 10047 17647 10053
rect 17589 10044 17601 10047
rect 17460 10016 17601 10044
rect 17460 10004 17466 10016
rect 17589 10013 17601 10016
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 16408 9976 16436 9992
rect 16408 9948 16712 9976
rect 16684 9917 16712 9948
rect 16117 9911 16175 9917
rect 16117 9908 16129 9911
rect 15948 9880 16129 9908
rect 16117 9877 16129 9880
rect 16163 9877 16175 9911
rect 16117 9871 16175 9877
rect 16669 9911 16727 9917
rect 16669 9877 16681 9911
rect 16715 9877 16727 9911
rect 17034 9908 17040 9920
rect 16995 9880 17040 9908
rect 16669 9871 16727 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 17129 9911 17187 9917
rect 17129 9877 17141 9911
rect 17175 9908 17187 9911
rect 17696 9908 17724 10084
rect 17862 10072 17868 10084
rect 17920 10112 17926 10124
rect 18414 10112 18420 10124
rect 17920 10084 18420 10112
rect 17920 10072 17926 10084
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 18046 10044 18052 10056
rect 18007 10016 18052 10044
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 17954 9936 17960 9988
rect 18012 9976 18018 9988
rect 18417 9979 18475 9985
rect 18417 9976 18429 9979
rect 18012 9948 18429 9976
rect 18012 9936 18018 9948
rect 18417 9945 18429 9948
rect 18463 9976 18475 9979
rect 18506 9976 18512 9988
rect 18463 9948 18512 9976
rect 18463 9945 18475 9948
rect 18417 9939 18475 9945
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 17175 9880 17724 9908
rect 17175 9877 17187 9880
rect 17129 9871 17187 9877
rect 17770 9868 17776 9920
rect 17828 9908 17834 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17828 9880 17877 9908
rect 17828 9868 17834 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 2225 9707 2283 9713
rect 2225 9673 2237 9707
rect 2271 9704 2283 9707
rect 2406 9704 2412 9716
rect 2271 9676 2412 9704
rect 2271 9673 2283 9676
rect 2225 9667 2283 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2556 9676 3188 9704
rect 2556 9664 2562 9676
rect 1673 9639 1731 9645
rect 1673 9605 1685 9639
rect 1719 9636 1731 9639
rect 2038 9636 2044 9648
rect 1719 9608 2044 9636
rect 1719 9605 1731 9608
rect 1673 9599 1731 9605
rect 2038 9596 2044 9608
rect 2096 9636 2102 9648
rect 2958 9636 2964 9648
rect 2096 9608 2964 9636
rect 2096 9596 2102 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3160 9636 3188 9676
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 3292 9676 4752 9704
rect 3292 9664 3298 9676
rect 3513 9639 3571 9645
rect 3160 9608 3464 9636
rect 1486 9568 1492 9580
rect 1399 9540 1492 9568
rect 1486 9528 1492 9540
rect 1544 9568 1550 9580
rect 2498 9568 2504 9580
rect 1544 9540 2504 9568
rect 1544 9528 1550 9540
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 2866 9568 2872 9580
rect 2779 9540 2872 9568
rect 2866 9528 2872 9540
rect 2924 9568 2930 9580
rect 3142 9568 3148 9580
rect 2924 9540 3148 9568
rect 2924 9528 2930 9540
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3436 9568 3464 9608
rect 3513 9605 3525 9639
rect 3559 9636 3571 9639
rect 4430 9636 4436 9648
rect 3559 9608 4436 9636
rect 3559 9605 3571 9608
rect 3513 9599 3571 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 4724 9636 4752 9676
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 5629 9707 5687 9713
rect 5629 9704 5641 9707
rect 4856 9676 5641 9704
rect 4856 9664 4862 9676
rect 5629 9673 5641 9676
rect 5675 9673 5687 9707
rect 5994 9704 6000 9716
rect 5629 9667 5687 9673
rect 5828 9676 6000 9704
rect 4982 9636 4988 9648
rect 4724 9608 4988 9636
rect 4982 9596 4988 9608
rect 5040 9636 5046 9648
rect 5537 9639 5595 9645
rect 5537 9636 5549 9639
rect 5040 9608 5549 9636
rect 5040 9596 5046 9608
rect 5537 9605 5549 9608
rect 5583 9605 5595 9639
rect 5828 9636 5856 9676
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6420 9676 6837 9704
rect 6420 9664 6426 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 8294 9704 8300 9716
rect 6825 9667 6883 9673
rect 6932 9676 8300 9704
rect 5537 9599 5595 9605
rect 5736 9608 5856 9636
rect 3970 9568 3976 9580
rect 3436 9540 3976 9568
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 4341 9571 4399 9577
rect 4341 9568 4353 9571
rect 4304 9540 4353 9568
rect 4304 9528 4310 9540
rect 4341 9537 4353 9540
rect 4387 9568 4399 9571
rect 5736 9568 5764 9608
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 5960 9608 6745 9636
rect 5960 9596 5966 9608
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6932 9636 6960 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8481 9707 8539 9713
rect 8481 9673 8493 9707
rect 8527 9704 8539 9707
rect 8938 9704 8944 9716
rect 8527 9676 8944 9704
rect 8527 9673 8539 9676
rect 8481 9667 8539 9673
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 9306 9704 9312 9716
rect 9267 9676 9312 9704
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10045 9707 10103 9713
rect 10045 9673 10057 9707
rect 10091 9704 10103 9707
rect 10226 9704 10232 9716
rect 10091 9676 10232 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10413 9707 10471 9713
rect 10413 9673 10425 9707
rect 10459 9704 10471 9707
rect 11238 9704 11244 9716
rect 10459 9676 11244 9704
rect 10459 9673 10471 9676
rect 10413 9667 10471 9673
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 11974 9704 11980 9716
rect 11935 9676 11980 9704
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 13136 9676 13185 9704
rect 13136 9664 13142 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 13173 9667 13231 9673
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 13906 9704 13912 9716
rect 13412 9676 13912 9704
rect 13412 9664 13418 9676
rect 13906 9664 13912 9676
rect 13964 9704 13970 9716
rect 14642 9704 14648 9716
rect 13964 9676 14648 9704
rect 13964 9664 13970 9676
rect 6733 9599 6791 9605
rect 6840 9608 6960 9636
rect 7024 9608 8524 9636
rect 4387 9540 5764 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 6638 9568 6644 9580
rect 5868 9540 6644 9568
rect 5868 9528 5874 9540
rect 6638 9528 6644 9540
rect 6696 9568 6702 9580
rect 6840 9568 6868 9608
rect 6696 9540 6868 9568
rect 6696 9528 6702 9540
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 1964 9432 1992 9463
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 2096 9472 2145 9500
rect 2096 9460 2102 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 2133 9463 2191 9469
rect 2746 9472 3617 9500
rect 2222 9432 2228 9444
rect 1964 9404 2228 9432
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2746 9432 2774 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 3145 9435 3203 9441
rect 3145 9432 3157 9435
rect 2639 9404 2774 9432
rect 2884 9404 3157 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2884 9364 2912 9404
rect 3145 9401 3157 9404
rect 3191 9401 3203 9435
rect 3145 9395 3203 9401
rect 2832 9336 2912 9364
rect 3053 9367 3111 9373
rect 2832 9324 2838 9336
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3510 9364 3516 9376
rect 3099 9336 3516 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3804 9364 3832 9463
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4120 9472 4445 9500
rect 4120 9460 4126 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 4798 9500 4804 9512
rect 4580 9472 4625 9500
rect 4759 9472 4804 9500
rect 4580 9460 4586 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 6178 9500 6184 9512
rect 5767 9472 6184 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6270 9460 6276 9512
rect 6328 9500 6334 9512
rect 6328 9472 6500 9500
rect 6328 9460 6334 9472
rect 3973 9435 4031 9441
rect 3973 9401 3985 9435
rect 4019 9432 4031 9435
rect 4154 9432 4160 9444
rect 4019 9404 4160 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 4396 9404 5948 9432
rect 4396 9392 4402 9404
rect 4890 9364 4896 9376
rect 3804 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5166 9364 5172 9376
rect 5127 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5920 9364 5948 9404
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 6089 9435 6147 9441
rect 6089 9432 6101 9435
rect 6052 9404 6101 9432
rect 6052 9392 6058 9404
rect 6089 9401 6101 9404
rect 6135 9401 6147 9435
rect 6362 9432 6368 9444
rect 6323 9404 6368 9432
rect 6089 9395 6147 9401
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 6472 9432 6500 9472
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6880 9472 6929 9500
rect 6880 9460 6886 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7024 9432 7052 9608
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 8018 9568 8024 9580
rect 7607 9540 8024 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8496 9568 8524 9608
rect 8570 9596 8576 9648
rect 8628 9636 8634 9648
rect 12802 9636 12808 9648
rect 8628 9608 9444 9636
rect 8628 9596 8634 9608
rect 9122 9568 9128 9580
rect 8496 9540 9128 9568
rect 8389 9531 8447 9537
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 7248 9472 7297 9500
rect 7248 9460 7254 9472
rect 7285 9469 7297 9472
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 8294 9500 8300 9512
rect 7515 9472 8300 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8404 9500 8432 9531
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9214 9528 9220 9580
rect 9272 9568 9278 9580
rect 9272 9540 9317 9568
rect 9272 9528 9278 9540
rect 8570 9500 8576 9512
rect 8404 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 8938 9500 8944 9512
rect 8711 9472 8944 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 9416 9509 9444 9608
rect 9784 9608 12808 9636
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9674 9500 9680 9512
rect 9447 9472 9680 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9784 9509 9812 9608
rect 12802 9596 12808 9608
rect 12860 9636 12866 9648
rect 12860 9608 13032 9636
rect 12860 9596 12866 9608
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9469 9827 9503
rect 9950 9500 9956 9512
rect 9911 9472 9956 9500
rect 9769 9463 9827 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9469 10563 9503
rect 10778 9500 10784 9512
rect 10739 9472 10784 9500
rect 10505 9463 10563 9469
rect 6472 9404 7052 9432
rect 7929 9435 7987 9441
rect 7929 9401 7941 9435
rect 7975 9432 7987 9435
rect 8110 9432 8116 9444
rect 7975 9404 8116 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 8202 9392 8208 9444
rect 8260 9432 8266 9444
rect 8849 9435 8907 9441
rect 8849 9432 8861 9435
rect 8260 9404 8861 9432
rect 8260 9392 8266 9404
rect 8849 9401 8861 9404
rect 8895 9401 8907 9435
rect 8849 9395 8907 9401
rect 9214 9392 9220 9444
rect 9272 9432 9278 9444
rect 10410 9432 10416 9444
rect 9272 9404 10416 9432
rect 9272 9392 9278 9404
rect 10410 9392 10416 9404
rect 10468 9432 10474 9444
rect 10520 9432 10548 9463
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 10468 9404 10548 9432
rect 11900 9432 11928 9531
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12492 9540 12725 9568
rect 12492 9528 12498 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 12066 9500 12072 9512
rect 12027 9472 12072 9500
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12802 9500 12808 9512
rect 12676 9472 12808 9500
rect 12676 9460 12682 9472
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 13004 9509 13032 9608
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13998 9636 14004 9648
rect 13688 9608 14004 9636
rect 13688 9596 13694 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 14292 9645 14320 9676
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 14737 9707 14795 9713
rect 14737 9673 14749 9707
rect 14783 9704 14795 9707
rect 15010 9704 15016 9716
rect 14783 9676 15016 9704
rect 14783 9673 14795 9676
rect 14737 9667 14795 9673
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 15197 9707 15255 9713
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15746 9704 15752 9716
rect 15243 9676 15752 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16390 9704 16396 9716
rect 16351 9676 16396 9704
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 18414 9704 18420 9716
rect 16540 9676 18000 9704
rect 18375 9676 18420 9704
rect 16540 9664 16546 9676
rect 14277 9639 14335 9645
rect 14277 9605 14289 9639
rect 14323 9605 14335 9639
rect 14277 9599 14335 9605
rect 14369 9639 14427 9645
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 14918 9636 14924 9648
rect 14415 9608 14924 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 15286 9636 15292 9648
rect 15247 9608 15292 9636
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 15712 9608 15945 9636
rect 15712 9596 15718 9608
rect 15933 9605 15945 9608
rect 15979 9605 15991 9639
rect 15933 9599 15991 9605
rect 16025 9639 16083 9645
rect 16025 9605 16037 9639
rect 16071 9636 16083 9639
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16071 9608 16957 9636
rect 16071 9605 16083 9608
rect 16025 9599 16083 9605
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 16945 9599 17003 9605
rect 17310 9596 17316 9648
rect 17368 9636 17374 9648
rect 17678 9636 17684 9648
rect 17368 9608 17684 9636
rect 17368 9596 17374 9608
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 13538 9568 13544 9580
rect 13499 9540 13544 9568
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 15194 9568 15200 9580
rect 14200 9540 15200 9568
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13078 9500 13084 9512
rect 13035 9472 13084 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13630 9500 13636 9512
rect 13591 9472 13636 9500
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 14200 9509 14228 9540
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 16850 9568 16856 9580
rect 16811 9540 16856 9568
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 16960 9540 17509 9568
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9469 14243 9503
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 14185 9463 14243 9469
rect 14476 9472 15393 9500
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 11900 9404 12357 9432
rect 10468 9392 10474 9404
rect 12345 9401 12357 9404
rect 12391 9401 12403 9435
rect 13740 9432 13768 9463
rect 14476 9432 14504 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 15562 9460 15568 9512
rect 15620 9500 15626 9512
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 15620 9472 15761 9500
rect 15620 9460 15626 9472
rect 15749 9469 15761 9472
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16960 9500 16988 9540
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 17972 9568 18000 9676
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 17972 9540 18337 9568
rect 17497 9531 17555 9537
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 16080 9472 16988 9500
rect 17221 9503 17279 9509
rect 16080 9460 16086 9472
rect 17221 9469 17233 9503
rect 17267 9500 17279 9503
rect 17954 9500 17960 9512
rect 17267 9472 17960 9500
rect 17267 9469 17279 9472
rect 17221 9463 17279 9469
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 12345 9395 12403 9401
rect 13096 9404 13768 9432
rect 14108 9404 14504 9432
rect 6454 9364 6460 9376
rect 5920 9336 6460 9364
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 8021 9367 8079 9373
rect 8021 9364 8033 9367
rect 6972 9336 8033 9364
rect 6972 9324 6978 9336
rect 8021 9333 8033 9336
rect 8067 9333 8079 9367
rect 8021 9327 8079 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10502 9364 10508 9376
rect 10192 9336 10508 9364
rect 10192 9324 10198 9336
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11422 9324 11428 9376
rect 11480 9364 11486 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11480 9336 11529 9364
rect 11480 9324 11486 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11517 9327 11575 9333
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 13096 9364 13124 9404
rect 11664 9336 13124 9364
rect 11664 9324 11670 9336
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 14108 9364 14136 9404
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 14608 9404 16681 9432
rect 14608 9392 14614 9404
rect 16669 9401 16681 9404
rect 16715 9401 16727 9435
rect 16669 9395 16727 9401
rect 17402 9392 17408 9444
rect 17460 9432 17466 9444
rect 17862 9432 17868 9444
rect 17460 9404 17868 9432
rect 17460 9392 17466 9404
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 18141 9435 18199 9441
rect 18141 9401 18153 9435
rect 18187 9432 18199 9435
rect 18598 9432 18604 9444
rect 18187 9404 18604 9432
rect 18187 9401 18199 9404
rect 18141 9395 18199 9401
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 13780 9336 14136 9364
rect 13780 9324 13786 9336
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14240 9336 14841 9364
rect 14240 9324 14246 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 18230 9364 18236 9376
rect 14976 9336 18236 9364
rect 14976 9324 14982 9336
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 3510 9160 3516 9172
rect 2280 9132 3516 9160
rect 2280 9120 2286 9132
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 8018 9160 8024 9172
rect 4264 9132 7880 9160
rect 7979 9132 8024 9160
rect 1673 9095 1731 9101
rect 1673 9061 1685 9095
rect 1719 9092 1731 9095
rect 3694 9092 3700 9104
rect 1719 9064 3700 9092
rect 1719 9061 1731 9064
rect 1673 9055 1731 9061
rect 3694 9052 3700 9064
rect 3752 9052 3758 9104
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 2406 9024 2412 9036
rect 1636 8996 2412 9024
rect 1636 8984 1642 8996
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 4264 9024 4292 9132
rect 4614 9052 4620 9104
rect 4672 9092 4678 9104
rect 6181 9095 6239 9101
rect 4672 9064 6132 9092
rect 4672 9052 4678 9064
rect 4430 9024 4436 9036
rect 3160 8996 4292 9024
rect 4391 8996 4436 9024
rect 1946 8916 1952 8968
rect 2004 8956 2010 8968
rect 2777 8959 2835 8965
rect 2777 8956 2789 8959
rect 2004 8928 2789 8956
rect 2004 8916 2010 8928
rect 2777 8925 2789 8928
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 1489 8891 1547 8897
rect 1489 8857 1501 8891
rect 1535 8888 1547 8891
rect 1578 8888 1584 8900
rect 1535 8860 1584 8888
rect 1535 8857 1547 8860
rect 1489 8851 1547 8857
rect 1578 8848 1584 8860
rect 1636 8888 1642 8900
rect 3160 8888 3188 8996
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4764 8996 5181 9024
rect 4764 8984 4770 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5626 9024 5632 9036
rect 5587 8996 5632 9024
rect 5169 8987 5227 8993
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 6104 9024 6132 9064
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 6454 9092 6460 9104
rect 6227 9064 6460 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 6454 9052 6460 9064
rect 6512 9052 6518 9104
rect 6104 8996 6684 9024
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3602 8956 3608 8968
rect 3283 8928 3608 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3602 8916 3608 8928
rect 3660 8956 3666 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 3660 8928 4997 8956
rect 3660 8916 3666 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 4985 8919 5043 8925
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 6546 8956 6552 8968
rect 6507 8928 6552 8956
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6656 8956 6684 8996
rect 7852 8956 7880 9132
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8352 9132 8953 9160
rect 8352 9120 8358 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 9766 9160 9772 9172
rect 9456 9132 9772 9160
rect 9456 9120 9462 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10008 9132 10885 9160
rect 10008 9120 10014 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 10873 9123 10931 9129
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 14550 9160 14556 9172
rect 11572 9132 14556 9160
rect 11572 9120 11578 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15194 9160 15200 9172
rect 14660 9132 15200 9160
rect 7929 9095 7987 9101
rect 7929 9061 7941 9095
rect 7975 9061 7987 9095
rect 7929 9055 7987 9061
rect 7944 9024 7972 9055
rect 9306 9052 9312 9104
rect 9364 9092 9370 9104
rect 9364 9064 9674 9092
rect 9364 9052 9370 9064
rect 8662 9024 8668 9036
rect 7944 8996 8668 9024
rect 8662 8984 8668 8996
rect 8720 9024 8726 9036
rect 9490 9024 9496 9036
rect 8720 8996 9496 9024
rect 8720 8984 8726 8996
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9646 9024 9674 9064
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 13630 9092 13636 9104
rect 12676 9064 13636 9092
rect 12676 9052 12682 9064
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 14458 9092 14464 9104
rect 14419 9064 14464 9092
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 9858 9024 9864 9036
rect 9646 8996 9864 9024
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10689 9027 10747 9033
rect 10100 8996 10640 9024
rect 10100 8984 10106 8996
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 6656 8928 7624 8956
rect 7852 8928 9413 8956
rect 1636 8860 3188 8888
rect 3513 8891 3571 8897
rect 1636 8848 1642 8860
rect 3513 8857 3525 8891
rect 3559 8888 3571 8891
rect 4157 8891 4215 8897
rect 4157 8888 4169 8891
rect 3559 8860 4169 8888
rect 3559 8857 3571 8860
rect 3513 8851 3571 8857
rect 4157 8857 4169 8860
rect 4203 8857 4215 8891
rect 4157 8851 4215 8857
rect 4890 8848 4896 8900
rect 4948 8888 4954 8900
rect 6822 8897 6828 8900
rect 6816 8888 6828 8897
rect 4948 8860 6684 8888
rect 6783 8860 6828 8888
rect 4948 8848 4954 8860
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8820 1826 8832
rect 2317 8823 2375 8829
rect 2317 8820 2329 8823
rect 1820 8792 2329 8820
rect 1820 8780 1826 8792
rect 2317 8789 2329 8792
rect 2363 8789 2375 8823
rect 2317 8783 2375 8789
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 2958 8820 2964 8832
rect 2464 8792 2509 8820
rect 2919 8792 2964 8820
rect 2464 8780 2470 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3292 8792 3801 8820
rect 3292 8780 3298 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 4120 8792 4261 8820
rect 4120 8780 4126 8792
rect 4249 8789 4261 8792
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 4488 8792 4629 8820
rect 4488 8780 4494 8792
rect 4617 8789 4629 8792
rect 4663 8789 4675 8823
rect 5074 8820 5080 8832
rect 5035 8792 5080 8820
rect 4617 8783 4675 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5718 8820 5724 8832
rect 5679 8792 5724 8820
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6273 8823 6331 8829
rect 6273 8820 6285 8823
rect 5960 8792 6285 8820
rect 5960 8780 5966 8792
rect 6273 8789 6285 8792
rect 6319 8789 6331 8823
rect 6656 8820 6684 8860
rect 6816 8851 6828 8860
rect 6822 8848 6828 8851
rect 6880 8848 6886 8900
rect 7596 8888 7624 8928
rect 9401 8925 9413 8928
rect 9447 8956 9459 8959
rect 9766 8956 9772 8968
rect 9447 8928 9772 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10192 8928 10517 8956
rect 10192 8916 10198 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10612 8956 10640 8996
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 11238 9024 11244 9036
rect 10735 8996 11244 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11514 9024 11520 9036
rect 11388 8996 11433 9024
rect 11475 8996 11520 9024
rect 11388 8984 11394 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 9024 12311 9027
rect 12434 9024 12440 9036
rect 12299 8996 12440 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 12434 8984 12440 8996
rect 12492 8984 12498 9036
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 12860 8996 13185 9024
rect 12860 8984 12866 8996
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13596 8996 14197 9024
rect 13596 8984 13602 8996
rect 14185 8993 14197 8996
rect 14231 9024 14243 9027
rect 14550 9024 14556 9036
rect 14231 8996 14556 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 14660 9033 14688 9132
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15286 9120 15292 9172
rect 15344 9160 15350 9172
rect 15381 9163 15439 9169
rect 15381 9160 15393 9163
rect 15344 9132 15393 9160
rect 15344 9120 15350 9132
rect 15381 9129 15393 9132
rect 15427 9129 15439 9163
rect 15381 9123 15439 9129
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 15804 9132 17448 9160
rect 15804 9120 15810 9132
rect 14918 9052 14924 9104
rect 14976 9092 14982 9104
rect 16942 9092 16948 9104
rect 14976 9064 16948 9092
rect 14976 9052 14982 9064
rect 16942 9052 16948 9064
rect 17000 9052 17006 9104
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 8993 14703 9027
rect 14826 9024 14832 9036
rect 14787 8996 14832 9024
rect 14645 8987 14703 8993
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15068 8996 15945 9024
rect 15068 8984 15074 8996
rect 15933 8993 15945 8996
rect 15979 9024 15991 9027
rect 16114 9024 16120 9036
rect 15979 8996 16120 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 16850 9024 16856 9036
rect 16356 8996 16712 9024
rect 16811 8996 16856 9024
rect 16356 8984 16362 8996
rect 13556 8956 13584 8984
rect 10612 8928 13584 8956
rect 10505 8919 10563 8925
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 13909 8959 13967 8965
rect 13688 8928 13733 8956
rect 13688 8916 13694 8928
rect 13909 8925 13921 8959
rect 13955 8956 13967 8959
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13955 8928 14289 8956
rect 13955 8925 13967 8928
rect 13909 8919 13967 8925
rect 14277 8925 14289 8928
rect 14323 8956 14335 8959
rect 15194 8956 15200 8968
rect 14323 8928 15200 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 15194 8916 15200 8928
rect 15252 8916 15258 8968
rect 16022 8956 16028 8968
rect 15304 8928 16028 8956
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 7596 8860 8493 8888
rect 8481 8857 8493 8860
rect 8527 8888 8539 8891
rect 9214 8888 9220 8900
rect 8527 8860 9220 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 9214 8848 9220 8860
rect 9272 8848 9278 8900
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 11241 8891 11299 8897
rect 11241 8888 11253 8891
rect 9364 8860 11253 8888
rect 9364 8848 9370 8860
rect 11241 8857 11253 8860
rect 11287 8888 11299 8891
rect 15304 8888 15332 8928
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16448 8928 16589 8956
rect 16448 8916 16454 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16684 8956 16712 8996
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 16942 8956 16948 8968
rect 16684 8928 16948 8956
rect 16577 8919 16635 8925
rect 16942 8916 16948 8928
rect 17000 8956 17006 8968
rect 17000 8928 17356 8956
rect 17000 8916 17006 8928
rect 11287 8860 15332 8888
rect 15841 8891 15899 8897
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 15841 8857 15853 8891
rect 15887 8888 15899 8891
rect 15887 8860 17080 8888
rect 15887 8857 15899 8860
rect 15841 8851 15899 8857
rect 7098 8820 7104 8832
rect 6656 8792 7104 8820
rect 6273 8783 6331 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8260 8792 8401 8820
rect 8260 8780 8266 8792
rect 8389 8789 8401 8792
rect 8435 8820 8447 8823
rect 9398 8820 9404 8832
rect 8435 8792 9404 8820
rect 8435 8789 8447 8792
rect 8389 8783 8447 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 10045 8823 10103 8829
rect 10045 8820 10057 8823
rect 9916 8792 10057 8820
rect 9916 8780 9922 8792
rect 10045 8789 10057 8792
rect 10091 8789 10103 8823
rect 10045 8783 10103 8789
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8820 10471 8823
rect 11422 8820 11428 8832
rect 10459 8792 11428 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12676 8792 13001 8820
rect 12676 8780 12682 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 12989 8783 13047 8789
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 14366 8820 14372 8832
rect 13587 8792 14372 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 14366 8780 14372 8792
rect 14424 8820 14430 8832
rect 14734 8820 14740 8832
rect 14424 8792 14740 8820
rect 14424 8780 14430 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 14918 8820 14924 8832
rect 14879 8792 14924 8820
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 15289 8823 15347 8829
rect 15289 8789 15301 8823
rect 15335 8820 15347 8823
rect 15378 8820 15384 8832
rect 15335 8792 15384 8820
rect 15335 8789 15347 8792
rect 15289 8783 15347 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16206 8820 16212 8832
rect 16167 8792 16212 8820
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17052 8829 17080 8860
rect 17037 8823 17095 8829
rect 16724 8792 16769 8820
rect 16724 8780 16730 8792
rect 17037 8789 17049 8823
rect 17083 8789 17095 8823
rect 17328 8820 17356 8928
rect 17420 8897 17448 9132
rect 17586 9024 17592 9036
rect 17547 8996 17592 9024
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 18046 8956 18052 8968
rect 18007 8928 18052 8956
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18230 8956 18236 8968
rect 18191 8928 18236 8956
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 17405 8891 17463 8897
rect 17405 8857 17417 8891
rect 17451 8888 17463 8891
rect 17954 8888 17960 8900
rect 17451 8860 17960 8888
rect 17451 8857 17463 8860
rect 17405 8851 17463 8857
rect 17954 8848 17960 8860
rect 18012 8888 18018 8900
rect 18322 8888 18328 8900
rect 18012 8860 18328 8888
rect 18012 8848 18018 8860
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 17497 8823 17555 8829
rect 17497 8820 17509 8823
rect 17328 8792 17509 8820
rect 17037 8783 17095 8789
rect 17497 8789 17509 8792
rect 17543 8789 17555 8823
rect 17862 8820 17868 8832
rect 17823 8792 17868 8820
rect 17497 8783 17555 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18417 8823 18475 8829
rect 18417 8789 18429 8823
rect 18463 8820 18475 8823
rect 18506 8820 18512 8832
rect 18463 8792 18512 8820
rect 18463 8789 18475 8792
rect 18417 8783 18475 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8585 2467 8619
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 2409 8579 2467 8585
rect 1486 8548 1492 8560
rect 1399 8520 1492 8548
rect 1486 8508 1492 8520
rect 1544 8548 1550 8560
rect 2424 8548 2452 8579
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 4430 8616 4436 8628
rect 3384 8588 3429 8616
rect 4391 8588 4436 8616
rect 3384 8576 3390 8588
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6822 8616 6828 8628
rect 6227 8588 6828 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8619 8588 10180 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 3881 8551 3939 8557
rect 1544 8520 2084 8548
rect 2424 8520 3188 8548
rect 1544 8508 1550 8520
rect 2056 8492 2084 8520
rect 1762 8480 1768 8492
rect 1723 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8440 1826 8492
rect 2038 8440 2044 8492
rect 2096 8440 2102 8492
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 3050 8480 3056 8492
rect 2547 8452 3056 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2280 8384 2697 8412
rect 2280 8372 2286 8384
rect 2685 8381 2697 8384
rect 2731 8412 2743 8415
rect 2958 8412 2964 8424
rect 2731 8384 2964 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 1946 8344 1952 8356
rect 1907 8316 1952 8344
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 3160 8344 3188 8520
rect 3881 8517 3893 8551
rect 3927 8548 3939 8551
rect 4154 8548 4160 8560
rect 3927 8520 4160 8548
rect 3927 8517 3939 8520
rect 3881 8511 3939 8517
rect 4154 8508 4160 8520
rect 4212 8508 4218 8560
rect 6546 8548 6552 8560
rect 4816 8520 6552 8548
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 4338 8480 4344 8492
rect 3568 8452 4200 8480
rect 4299 8452 4344 8480
rect 3568 8440 3574 8452
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 3476 8384 3521 8412
rect 3476 8372 3482 8384
rect 2464 8316 3188 8344
rect 2464 8304 2470 8316
rect 3878 8304 3884 8356
rect 3936 8344 3942 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 3936 8316 3985 8344
rect 3936 8304 3942 8316
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 2869 8279 2927 8285
rect 2869 8245 2881 8279
rect 2915 8276 2927 8279
rect 3510 8276 3516 8288
rect 2915 8248 3516 8276
rect 2915 8245 2927 8248
rect 2869 8239 2927 8245
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 4172 8276 4200 8452
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4816 8489 4844 8520
rect 6546 8508 6552 8520
rect 6604 8548 6610 8560
rect 8846 8548 8852 8560
rect 6604 8520 8852 8548
rect 6604 8508 6610 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 5068 8483 5126 8489
rect 5068 8449 5080 8483
rect 5114 8480 5126 8483
rect 6086 8480 6092 8492
rect 5114 8452 6092 8480
rect 5114 8449 5126 8452
rect 5068 8443 5126 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 7208 8489 7236 8520
rect 8846 8508 8852 8520
rect 8904 8548 8910 8560
rect 10152 8548 10180 8588
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 10284 8588 10517 8616
rect 10284 8576 10290 8588
rect 10505 8585 10517 8588
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13354 8616 13360 8628
rect 12492 8588 13360 8616
rect 12492 8576 12498 8588
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 13780 8588 14841 8616
rect 13780 8576 13786 8588
rect 14829 8585 14841 8588
rect 14875 8616 14887 8619
rect 15378 8616 15384 8628
rect 14875 8588 15384 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 15712 8588 16405 8616
rect 15712 8576 15718 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16666 8616 16672 8628
rect 16627 8588 16672 8616
rect 16393 8579 16451 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 17034 8576 17040 8628
rect 17092 8576 17098 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17184 8588 17509 8616
rect 17184 8576 17190 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 17736 8588 17969 8616
rect 17736 8576 17742 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 11146 8548 11152 8560
rect 8904 8520 9168 8548
rect 10152 8520 11152 8548
rect 8904 8508 8910 8520
rect 7466 8489 7472 8492
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6564 8452 6745 8480
rect 4522 8412 4528 8424
rect 4483 8384 4528 8412
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6564 8412 6592 8452
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 7460 8480 7472 8489
rect 7427 8452 7472 8480
rect 7193 8443 7251 8449
rect 7460 8443 7472 8452
rect 7466 8440 7472 8443
rect 7524 8440 7530 8492
rect 9140 8489 9168 8520
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 15188 8551 15246 8557
rect 15188 8548 15200 8551
rect 11624 8520 14964 8548
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9381 8483 9439 8489
rect 9381 8480 9393 8483
rect 9272 8452 9393 8480
rect 9272 8440 9278 8452
rect 9381 8449 9393 8452
rect 9427 8449 9439 8483
rect 9381 8443 9439 8449
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 11624 8489 11652 8520
rect 13464 8489 13492 8520
rect 11609 8483 11667 8489
rect 11609 8480 11621 8483
rect 11388 8452 11621 8480
rect 11388 8440 11394 8452
rect 11609 8449 11621 8452
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 11876 8483 11934 8489
rect 11876 8449 11888 8483
rect 11922 8480 11934 8483
rect 13449 8483 13507 8489
rect 11922 8452 13400 8480
rect 11922 8449 11934 8452
rect 11876 8443 11934 8449
rect 5960 8384 6592 8412
rect 5960 8372 5966 8384
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6696 8384 6837 8412
rect 6696 8372 6702 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 13372 8412 13400 8452
rect 13449 8449 13461 8483
rect 13495 8449 13507 8483
rect 13449 8443 13507 8449
rect 13716 8483 13774 8489
rect 13716 8449 13728 8483
rect 13762 8480 13774 8483
rect 14826 8480 14832 8492
rect 13762 8452 14832 8480
rect 13762 8449 13774 8452
rect 13716 8443 13774 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 14936 8489 14964 8520
rect 15028 8520 15200 8548
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 13372 8384 13492 8412
rect 6917 8375 6975 8381
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 5868 8316 6377 8344
rect 5868 8304 5874 8316
rect 6365 8313 6377 8316
rect 6411 8313 6423 8347
rect 6932 8344 6960 8375
rect 8757 8347 8815 8353
rect 6365 8307 6423 8313
rect 6472 8316 7236 8344
rect 5902 8276 5908 8288
rect 4172 8248 5908 8276
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6472 8276 6500 8316
rect 6236 8248 6500 8276
rect 7208 8276 7236 8316
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9030 8344 9036 8356
rect 8803 8316 9036 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 12986 8344 12992 8356
rect 12768 8316 12992 8344
rect 12768 8304 12774 8316
rect 12986 8304 12992 8316
rect 13044 8304 13050 8356
rect 13170 8344 13176 8356
rect 13131 8316 13176 8344
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 7926 8276 7932 8288
rect 7208 8248 7932 8276
rect 6236 8236 6242 8248
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9398 8276 9404 8288
rect 8987 8248 9404 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 13464 8276 13492 8384
rect 14458 8372 14464 8424
rect 14516 8412 14522 8424
rect 15028 8412 15056 8520
rect 15188 8517 15200 8520
rect 15234 8548 15246 8551
rect 15286 8548 15292 8560
rect 15234 8520 15292 8548
rect 15234 8517 15246 8520
rect 15188 8511 15246 8517
rect 15286 8508 15292 8520
rect 15344 8508 15350 8560
rect 15562 8508 15568 8560
rect 15620 8548 15626 8560
rect 17052 8548 17080 8576
rect 17865 8551 17923 8557
rect 17865 8548 17877 8551
rect 15620 8520 16068 8548
rect 17052 8520 17877 8548
rect 15620 8508 15626 8520
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15528 8452 15976 8480
rect 15528 8440 15534 8452
rect 14516 8384 15056 8412
rect 14516 8372 14522 8384
rect 15948 8356 15976 8452
rect 16040 8412 16068 8520
rect 17865 8517 17877 8520
rect 17911 8517 17923 8551
rect 17865 8511 17923 8517
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 16816 8452 17049 8480
rect 16816 8440 16822 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17494 8480 17500 8492
rect 17175 8452 17500 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18012 8452 18521 8480
rect 18012 8440 18018 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16040 8384 17233 8412
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17221 8375 17279 8381
rect 17328 8384 18061 8412
rect 15930 8304 15936 8356
rect 15988 8344 15994 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 15988 8316 16313 8344
rect 15988 8304 15994 8316
rect 16301 8313 16313 8316
rect 16347 8313 16359 8347
rect 16301 8307 16359 8313
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 17328 8344 17356 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18874 8412 18880 8424
rect 18049 8375 18107 8381
rect 18156 8384 18880 8412
rect 16448 8316 17356 8344
rect 16448 8304 16454 8316
rect 17494 8304 17500 8356
rect 17552 8344 17558 8356
rect 18156 8344 18184 8384
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 17552 8316 18184 8344
rect 18325 8347 18383 8353
rect 17552 8304 17558 8316
rect 18325 8313 18337 8347
rect 18371 8344 18383 8347
rect 18782 8344 18788 8356
rect 18371 8316 18788 8344
rect 18371 8313 18383 8316
rect 18325 8307 18383 8313
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 15102 8276 15108 8288
rect 13464 8248 15108 8276
rect 15102 8236 15108 8248
rect 15160 8276 15166 8288
rect 15654 8276 15660 8288
rect 15160 8248 15660 8276
rect 15160 8236 15166 8248
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2958 8072 2964 8084
rect 2871 8044 2964 8072
rect 2958 8032 2964 8044
rect 3016 8072 3022 8084
rect 3016 8044 4292 8072
rect 3016 8032 3022 8044
rect 2409 8007 2467 8013
rect 2409 7973 2421 8007
rect 2455 7973 2467 8007
rect 4154 8004 4160 8016
rect 2409 7967 2467 7973
rect 3620 7976 4160 8004
rect 2424 7936 2452 7967
rect 3326 7936 3332 7948
rect 1688 7908 2452 7936
rect 2608 7908 3332 7936
rect 1688 7877 1716 7908
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2130 7868 2136 7880
rect 2087 7840 2136 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2608 7877 2636 7908
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3620 7877 3648 7976
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 4264 8004 4292 8044
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4396 8044 4721 8072
rect 4396 8032 4402 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 4709 8035 4767 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5718 8072 5724 8084
rect 5583 8044 5724 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 7285 8075 7343 8081
rect 5960 8044 6960 8072
rect 5960 8032 5966 8044
rect 4264 7976 5304 8004
rect 3786 7936 3792 7948
rect 3747 7908 3792 7936
rect 3786 7896 3792 7908
rect 3844 7896 3850 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4246 7936 4252 7948
rect 4111 7908 4252 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4246 7896 4252 7908
rect 4304 7936 4310 7948
rect 4706 7936 4712 7948
rect 4304 7908 4712 7936
rect 4304 7896 4310 7908
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7905 5043 7939
rect 4985 7899 5043 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5166 7936 5172 7948
rect 5123 7908 5172 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4798 7868 4804 7880
rect 4387 7840 4804 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5000 7868 5028 7899
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5276 7936 5304 7976
rect 6932 7936 6960 8044
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7374 8072 7380 8084
rect 7331 8044 7380 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 7484 8044 9597 8072
rect 7098 7964 7104 8016
rect 7156 8004 7162 8016
rect 7484 8004 7512 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 15470 8072 15476 8084
rect 9585 8035 9643 8041
rect 9692 8044 15476 8072
rect 7156 7976 7512 8004
rect 7156 7964 7162 7976
rect 9030 7964 9036 8016
rect 9088 8004 9094 8016
rect 9692 8004 9720 8044
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 15804 8044 17049 8072
rect 15804 8032 15810 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 17494 8072 17500 8084
rect 17368 8044 17500 8072
rect 17368 8032 17374 8044
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 18414 8072 18420 8084
rect 18375 8044 18420 8072
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 9088 7976 9720 8004
rect 12713 8007 12771 8013
rect 9088 7964 9094 7976
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 14458 8004 14464 8016
rect 12759 7976 14464 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 16945 8007 17003 8013
rect 16945 7973 16957 8007
rect 16991 7973 17003 8007
rect 16945 7967 17003 7973
rect 7558 7936 7564 7948
rect 5276 7908 6040 7936
rect 6932 7908 7564 7936
rect 5258 7868 5264 7880
rect 5000 7840 5264 7868
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6012 7868 6040 7908
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 10965 7939 11023 7945
rect 8680 7908 9996 7936
rect 8680 7868 8708 7908
rect 6012 7840 8708 7868
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8846 7868 8852 7880
rect 8803 7840 8852 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9968 7868 9996 7908
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11330 7936 11336 7948
rect 11011 7908 11336 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 10410 7868 10416 7880
rect 9968 7840 10416 7868
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11422 7868 11428 7880
rect 11296 7840 11428 7868
rect 11296 7828 11302 7840
rect 11422 7828 11428 7840
rect 11480 7868 11486 7880
rect 11589 7871 11647 7877
rect 11589 7868 11601 7871
rect 11480 7840 11601 7868
rect 11480 7828 11486 7840
rect 11589 7837 11601 7840
rect 11635 7837 11647 7871
rect 13630 7868 13636 7880
rect 13591 7840 13636 7868
rect 11589 7831 11647 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 15120 7840 15485 7868
rect 15120 7812 15148 7840
rect 15473 7837 15485 7840
rect 15519 7868 15531 7871
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15519 7840 15577 7868
rect 15519 7837 15531 7840
rect 15473 7831 15531 7837
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 16960 7868 16988 7967
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 17586 7936 17592 7948
rect 17368 7908 17592 7936
rect 17368 7896 17374 7908
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 17402 7868 17408 7880
rect 15712 7840 16988 7868
rect 17363 7840 17408 7868
rect 15712 7828 15718 7840
rect 17402 7828 17408 7840
rect 17460 7868 17466 7880
rect 17678 7868 17684 7880
rect 17460 7840 17684 7868
rect 17460 7828 17466 7840
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17862 7868 17868 7880
rect 17823 7840 17868 7868
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18322 7868 18328 7880
rect 18279 7840 18328 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 3142 7800 3148 7812
rect 2823 7772 3148 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 3142 7760 3148 7772
rect 3200 7760 3206 7812
rect 3326 7760 3332 7812
rect 3384 7800 3390 7812
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 3384 7772 4261 7800
rect 3384 7760 3390 7772
rect 4249 7769 4261 7772
rect 4295 7800 4307 7803
rect 4430 7800 4436 7812
rect 4295 7772 4436 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 5169 7803 5227 7809
rect 5169 7769 5181 7803
rect 5215 7800 5227 7803
rect 5810 7800 5816 7812
rect 5215 7772 5816 7800
rect 5215 7769 5227 7772
rect 5169 7763 5227 7769
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 6172 7803 6230 7809
rect 6172 7769 6184 7803
rect 6218 7800 6230 7803
rect 7006 7800 7012 7812
rect 6218 7772 7012 7800
rect 6218 7769 6230 7772
rect 6172 7763 6230 7769
rect 7006 7760 7012 7772
rect 7064 7760 7070 7812
rect 8512 7803 8570 7809
rect 8512 7769 8524 7803
rect 8558 7800 8570 7803
rect 10226 7800 10232 7812
rect 8558 7772 10232 7800
rect 8558 7769 8570 7772
rect 8512 7763 8570 7769
rect 10226 7760 10232 7772
rect 10284 7800 10290 7812
rect 10594 7800 10600 7812
rect 10284 7772 10600 7800
rect 10284 7760 10290 7772
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 10720 7803 10778 7809
rect 10720 7769 10732 7803
rect 10766 7800 10778 7803
rect 13909 7803 13967 7809
rect 10766 7772 11192 7800
rect 10766 7769 10778 7772
rect 10720 7763 10778 7769
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2038 7692 2044 7744
rect 2096 7732 2102 7744
rect 2133 7735 2191 7741
rect 2133 7732 2145 7735
rect 2096 7704 2145 7732
rect 2096 7692 2102 7704
rect 2133 7701 2145 7704
rect 2179 7701 2191 7735
rect 2133 7695 2191 7701
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 3053 7735 3111 7741
rect 3053 7732 3065 7735
rect 2556 7704 3065 7732
rect 2556 7692 2562 7704
rect 3053 7701 3065 7704
rect 3099 7701 3111 7735
rect 3418 7732 3424 7744
rect 3379 7704 3424 7732
rect 3053 7695 3111 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 7374 7732 7380 7744
rect 7335 7704 7380 7732
rect 7374 7692 7380 7704
rect 7432 7732 7438 7744
rect 8754 7732 8760 7744
rect 7432 7704 8760 7732
rect 7432 7692 7438 7704
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 11164 7741 11192 7772
rect 13909 7769 13921 7803
rect 13955 7800 13967 7803
rect 13955 7772 15056 7800
rect 13955 7769 13967 7772
rect 13909 7763 13967 7769
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11238 7732 11244 7744
rect 11195 7704 11244 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 14056 7704 14105 7732
rect 14056 7692 14062 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 15028 7732 15056 7772
rect 15102 7760 15108 7812
rect 15160 7760 15166 7812
rect 15194 7760 15200 7812
rect 15252 7809 15258 7812
rect 15252 7800 15264 7809
rect 15832 7803 15890 7809
rect 15252 7772 15297 7800
rect 15252 7763 15264 7772
rect 15832 7769 15844 7803
rect 15878 7800 15890 7803
rect 15930 7800 15936 7812
rect 15878 7772 15936 7800
rect 15878 7769 15890 7772
rect 15832 7763 15890 7769
rect 15252 7760 15258 7763
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 16022 7760 16028 7812
rect 16080 7800 16086 7812
rect 16080 7772 18276 7800
rect 16080 7760 16086 7772
rect 18248 7744 18276 7772
rect 16390 7732 16396 7744
rect 15028 7704 16396 7732
rect 14093 7695 14151 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 17862 7732 17868 7744
rect 17552 7704 17868 7732
rect 17552 7692 17558 7704
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 18046 7732 18052 7744
rect 18007 7704 18052 7732
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 18230 7692 18236 7744
rect 18288 7692 18294 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 2961 7531 3019 7537
rect 2961 7528 2973 7531
rect 2924 7500 2973 7528
rect 2924 7488 2930 7500
rect 2961 7497 2973 7500
rect 3007 7497 3019 7531
rect 2961 7491 3019 7497
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 3375 7500 5089 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 7929 7531 7987 7537
rect 5316 7500 7052 7528
rect 5316 7488 5322 7500
rect 1946 7420 1952 7472
rect 2004 7460 2010 7472
rect 2041 7463 2099 7469
rect 2041 7460 2053 7463
rect 2004 7432 2053 7460
rect 2004 7420 2010 7432
rect 2041 7429 2053 7432
rect 2087 7460 2099 7463
rect 2222 7460 2228 7472
rect 2087 7432 2228 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 2648 7432 3556 7460
rect 2648 7420 2654 7432
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 3418 7392 3424 7404
rect 3016 7364 3424 7392
rect 3016 7352 3022 7364
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 2866 7324 2872 7336
rect 2731 7296 2765 7324
rect 2827 7296 2872 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 1486 7256 1492 7268
rect 1447 7228 1492 7256
rect 1486 7216 1492 7228
rect 1544 7216 1550 7268
rect 1964 7256 1992 7287
rect 2700 7256 2728 7287
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3108 7296 3464 7324
rect 3108 7284 3114 7296
rect 3436 7265 3464 7296
rect 3421 7259 3479 7265
rect 1964 7228 2774 7256
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7188 2559 7191
rect 2590 7188 2596 7200
rect 2547 7160 2596 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 2746 7188 2774 7228
rect 3421 7225 3433 7259
rect 3467 7225 3479 7259
rect 3421 7219 3479 7225
rect 3142 7188 3148 7200
rect 2746 7160 3148 7188
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3528 7188 3556 7432
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 4433 7463 4491 7469
rect 4433 7460 4445 7463
rect 3660 7432 4445 7460
rect 3660 7420 3666 7432
rect 4433 7429 4445 7432
rect 4479 7429 4491 7463
rect 4433 7423 4491 7429
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 6914 7460 6920 7472
rect 5031 7432 6920 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7024 7460 7052 7500
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8478 7528 8484 7540
rect 7975 7500 8484 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 12894 7528 12900 7540
rect 8588 7500 12900 7528
rect 8588 7460 8616 7500
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13725 7531 13783 7537
rect 13725 7497 13737 7531
rect 13771 7528 13783 7531
rect 13814 7528 13820 7540
rect 13771 7500 13820 7528
rect 13771 7497 13783 7500
rect 13725 7491 13783 7497
rect 13814 7488 13820 7500
rect 13872 7488 13878 7540
rect 15381 7531 15439 7537
rect 15381 7497 15393 7531
rect 15427 7528 15439 7531
rect 16022 7528 16028 7540
rect 15427 7500 16028 7528
rect 15427 7497 15439 7500
rect 15381 7491 15439 7497
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16255 7500 16681 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16816 7500 17049 7528
rect 16816 7488 16822 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17957 7531 18015 7537
rect 17957 7528 17969 7531
rect 17184 7500 17969 7528
rect 17184 7488 17190 7500
rect 17957 7497 17969 7500
rect 18003 7497 18015 7531
rect 18322 7528 18328 7540
rect 18283 7500 18328 7528
rect 17957 7491 18015 7497
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 7024 7432 8616 7460
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 13081 7463 13139 7469
rect 8904 7432 11376 7460
rect 8904 7420 8910 7432
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 4154 7392 4160 7404
rect 3835 7364 4160 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 4338 7352 4344 7364
rect 4396 7392 4402 7404
rect 5534 7392 5540 7404
rect 4396 7364 5396 7392
rect 5495 7364 5540 7392
rect 4396 7352 4402 7364
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3752 7296 3893 7324
rect 3752 7284 3758 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4706 7324 4712 7336
rect 4019 7296 4712 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 3896 7256 3924 7287
rect 4062 7256 4068 7268
rect 3896 7228 4068 7256
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 4172 7188 4200 7296
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5166 7324 5172 7336
rect 5127 7296 5172 7324
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5368 7324 5396 7364
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 6638 7392 6644 7404
rect 6472 7364 6644 7392
rect 6472 7324 6500 7364
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 6816 7395 6874 7401
rect 6816 7361 6828 7395
rect 6862 7392 6874 7395
rect 7374 7392 7380 7404
rect 6862 7364 7380 7392
rect 6862 7361 6874 7364
rect 6816 7355 6874 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 9140 7401 9168 7432
rect 11348 7404 11376 7432
rect 13081 7429 13093 7463
rect 13127 7460 13139 7463
rect 17586 7460 17592 7472
rect 13127 7432 17592 7460
rect 13127 7429 13139 7432
rect 13081 7423 13139 7429
rect 17586 7420 17592 7432
rect 17644 7460 17650 7472
rect 17644 7432 18552 7460
rect 17644 7420 17650 7432
rect 9398 7401 9404 7404
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9392 7392 9404 7401
rect 9359 7364 9404 7392
rect 9125 7355 9183 7361
rect 9392 7355 9404 7364
rect 9398 7352 9404 7355
rect 9456 7352 9462 7404
rect 11330 7352 11336 7404
rect 11388 7392 11394 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11388 7364 11529 7392
rect 11388 7352 11394 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11773 7395 11831 7401
rect 11773 7392 11785 7395
rect 11664 7364 11785 7392
rect 11664 7352 11670 7364
rect 11773 7361 11785 7364
rect 11819 7361 11831 7395
rect 11773 7355 11831 7361
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 14838 7395 14896 7401
rect 14838 7392 14850 7395
rect 14148 7364 14850 7392
rect 14148 7352 14154 7364
rect 14838 7361 14850 7364
rect 14884 7361 14896 7395
rect 15102 7392 15108 7404
rect 15063 7364 15108 7392
rect 14838 7355 14896 7361
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15470 7392 15476 7404
rect 15431 7364 15476 7392
rect 15197 7355 15255 7361
rect 5368 7296 6500 7324
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 6564 7256 6592 7287
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13265 7327 13323 7333
rect 13265 7324 13277 7327
rect 13044 7296 13277 7324
rect 13044 7284 13050 7296
rect 13265 7293 13277 7296
rect 13311 7324 13323 7327
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 13311 7296 13461 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 13449 7293 13461 7296
rect 13495 7324 13507 7327
rect 13538 7324 13544 7336
rect 13495 7296 13544 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 5960 7228 6592 7256
rect 5960 7216 5966 7228
rect 4614 7188 4620 7200
rect 3528 7160 4200 7188
rect 4575 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 6564 7188 6592 7228
rect 10505 7259 10563 7265
rect 10505 7225 10517 7259
rect 10551 7256 10563 7259
rect 10686 7256 10692 7268
rect 10551 7228 10692 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 15212 7256 15240 7355
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 18524 7401 18552 7432
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 16408 7364 17877 7392
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 16080 7296 16313 7324
rect 16080 7284 16086 7296
rect 16301 7293 16313 7296
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 16408 7256 16436 7364
rect 17865 7361 17877 7364
rect 17911 7392 17923 7395
rect 18509 7395 18567 7401
rect 17911 7364 18184 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 17586 7324 17592 7336
rect 17359 7296 17592 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18156 7324 18184 7364
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 19058 7324 19064 7336
rect 18156 7296 19064 7324
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 15212 7228 16436 7256
rect 6822 7188 6828 7200
rect 6564 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 11238 7188 11244 7200
rect 7616 7160 11244 7188
rect 7616 7148 7622 7160
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 13446 7148 13452 7200
rect 13504 7188 13510 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13504 7160 13645 7188
rect 13504 7148 13510 7160
rect 13633 7157 13645 7160
rect 13679 7188 13691 7191
rect 15212 7188 15240 7228
rect 17402 7216 17408 7268
rect 17460 7256 17466 7268
rect 17460 7228 17540 7256
rect 17460 7216 17466 7228
rect 15654 7188 15660 7200
rect 13679 7160 15240 7188
rect 15615 7160 15660 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 17512 7197 17540 7228
rect 17497 7191 17555 7197
rect 15804 7160 15849 7188
rect 15804 7148 15810 7160
rect 17497 7157 17509 7191
rect 17543 7157 17555 7191
rect 17497 7151 17555 7157
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 2593 6987 2651 6993
rect 2593 6984 2605 6987
rect 1728 6956 2605 6984
rect 1728 6944 1734 6956
rect 2593 6953 2605 6956
rect 2639 6953 2651 6987
rect 2593 6947 2651 6953
rect 3804 6956 6960 6984
rect 1486 6916 1492 6928
rect 1447 6888 1492 6916
rect 1486 6876 1492 6888
rect 1544 6876 1550 6928
rect 2222 6916 2228 6928
rect 2183 6888 2228 6916
rect 2222 6876 2228 6888
rect 2280 6876 2286 6928
rect 3050 6916 3056 6928
rect 2963 6888 3056 6916
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2976 6857 3004 6888
rect 3050 6876 3056 6888
rect 3108 6916 3114 6928
rect 3804 6916 3832 6956
rect 3108 6888 3832 6916
rect 3108 6876 3114 6888
rect 3970 6876 3976 6928
rect 4028 6876 4034 6928
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2188 6820 2329 6848
rect 2188 6808 2194 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3694 6848 3700 6860
rect 3292 6820 3700 6848
rect 3292 6808 3298 6820
rect 3694 6808 3700 6820
rect 3752 6848 3758 6860
rect 3988 6848 4016 6876
rect 3752 6820 4016 6848
rect 6932 6848 6960 6956
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7064 6956 7297 6984
rect 7064 6944 7070 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10226 6984 10232 6996
rect 9999 6956 10232 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 11422 6984 11428 6996
rect 11383 6956 11428 6984
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 14826 6984 14832 6996
rect 13289 6956 14832 6984
rect 8757 6851 8815 6857
rect 6932 6820 7512 6848
rect 3752 6808 3758 6820
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1762 6780 1768 6792
rect 1719 6752 1768 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3050 6780 3056 6792
rect 2823 6752 3056 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4430 6780 4436 6792
rect 4391 6752 4436 6780
rect 4430 6740 4436 6752
rect 4488 6780 4494 6792
rect 5902 6780 5908 6792
rect 4488 6752 5908 6780
rect 4488 6740 4494 6752
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 3142 6712 3148 6724
rect 3055 6684 3148 6712
rect 3142 6672 3148 6684
rect 3200 6712 3206 6724
rect 3200 6684 4108 6712
rect 3200 6672 3206 6684
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3326 6644 3332 6656
rect 3283 6616 3332 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3602 6644 3608 6656
rect 3563 6616 3608 6644
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4080 6653 4108 6684
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 4212 6684 4261 6712
rect 4212 6672 4218 6684
rect 4249 6681 4261 6684
rect 4295 6712 4307 6715
rect 4338 6712 4344 6724
rect 4295 6684 4344 6712
rect 4295 6681 4307 6684
rect 4249 6675 4307 6681
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4700 6715 4758 6721
rect 4700 6681 4712 6715
rect 4746 6712 4758 6715
rect 5258 6712 5264 6724
rect 4746 6684 5264 6712
rect 4746 6681 4758 6684
rect 4700 6675 4758 6681
rect 5258 6672 5264 6684
rect 5316 6672 5322 6724
rect 6172 6715 6230 6721
rect 6172 6681 6184 6715
rect 6218 6712 6230 6715
rect 6218 6684 6776 6712
rect 6218 6681 6230 6684
rect 6172 6675 6230 6681
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 5718 6644 5724 6656
rect 4111 6616 5724 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 6270 6644 6276 6656
rect 5859 6616 6276 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6748 6644 6776 6684
rect 7190 6644 7196 6656
rect 6748 6616 7196 6644
rect 7190 6604 7196 6616
rect 7248 6644 7254 6656
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 7248 6616 7389 6644
rect 7248 6604 7254 6616
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 7484 6644 7512 6820
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 8846 6848 8852 6860
rect 8803 6820 8852 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 11330 6848 11336 6860
rect 11291 6820 11336 6848
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 12986 6848 12992 6860
rect 12947 6820 12992 6848
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 8501 6783 8559 6789
rect 8501 6749 8513 6783
rect 8547 6780 8559 6783
rect 8662 6780 8668 6792
rect 8547 6752 8668 6780
rect 8547 6749 8559 6752
rect 8501 6743 8559 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 11066 6783 11124 6789
rect 11066 6749 11078 6783
rect 11112 6780 11124 6783
rect 11348 6780 11376 6808
rect 12805 6783 12863 6789
rect 12805 6780 12817 6783
rect 11112 6752 11192 6780
rect 11348 6752 12817 6780
rect 11112 6749 11124 6752
rect 11066 6743 11124 6749
rect 11164 6724 11192 6752
rect 12805 6749 12817 6752
rect 12851 6749 12863 6783
rect 13289 6780 13317 6956
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15160 6956 15516 6984
rect 15160 6944 15166 6956
rect 13357 6919 13415 6925
rect 13357 6885 13369 6919
rect 13403 6916 13415 6919
rect 13722 6916 13728 6928
rect 13403 6888 13728 6916
rect 13403 6885 13415 6888
rect 13357 6879 13415 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 15488 6857 15516 6956
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 17310 6984 17316 6996
rect 15988 6956 17316 6984
rect 15988 6944 15994 6956
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 18414 6984 18420 6996
rect 18375 6956 18420 6984
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 17034 6876 17040 6928
rect 17092 6916 17098 6928
rect 18598 6916 18604 6928
rect 17092 6888 18604 6916
rect 17092 6876 17098 6888
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6848 15531 6851
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15519 6820 15577 6848
rect 15519 6817 15531 6820
rect 15473 6811 15531 6817
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 17586 6848 17592 6860
rect 17547 6820 17592 6848
rect 15565 6811 15623 6817
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 18046 6848 18052 6860
rect 17828 6820 18052 6848
rect 17828 6808 17834 6820
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 12805 6743 12863 6749
rect 12912 6752 13317 6780
rect 13372 6752 13461 6780
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 9214 6712 9220 6724
rect 8352 6684 9220 6712
rect 8352 6672 8358 6684
rect 9214 6672 9220 6684
rect 9272 6672 9278 6724
rect 11146 6672 11152 6724
rect 11204 6672 11210 6724
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 12538 6715 12596 6721
rect 12538 6712 12550 6715
rect 12032 6684 12550 6712
rect 12032 6672 12038 6684
rect 12538 6681 12550 6684
rect 12584 6681 12596 6715
rect 12538 6675 12596 6681
rect 12912 6656 12940 6752
rect 13372 6656 13400 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13722 6780 13728 6792
rect 13635 6752 13728 6780
rect 13449 6743 13507 6749
rect 13722 6740 13728 6752
rect 13780 6780 13786 6792
rect 14182 6780 14188 6792
rect 13780 6752 14188 6780
rect 13780 6740 13786 6752
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 15217 6783 15275 6789
rect 15217 6749 15229 6783
rect 15263 6780 15275 6783
rect 15378 6780 15384 6792
rect 15263 6752 15384 6780
rect 15263 6749 15275 6752
rect 15217 6743 15275 6749
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 16724 6752 17509 6780
rect 16724 6740 16730 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6780 17923 6783
rect 17954 6780 17960 6792
rect 17911 6752 17960 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 14826 6712 14832 6724
rect 13924 6684 14832 6712
rect 8938 6644 8944 6656
rect 7484 6616 8944 6644
rect 7377 6607 7435 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 12894 6644 12900 6656
rect 10836 6616 12900 6644
rect 10836 6604 10842 6616
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13173 6647 13231 6653
rect 13173 6613 13185 6647
rect 13219 6644 13231 6647
rect 13354 6644 13360 6656
rect 13219 6616 13360 6644
rect 13219 6613 13231 6616
rect 13173 6607 13231 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13630 6644 13636 6656
rect 13591 6616 13636 6644
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 13924 6653 13952 6684
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 15810 6715 15868 6721
rect 15810 6712 15822 6715
rect 15120 6684 15822 6712
rect 13909 6647 13967 6653
rect 13909 6613 13921 6647
rect 13955 6613 13967 6647
rect 13909 6607 13967 6613
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6644 14151 6647
rect 14274 6644 14280 6656
rect 14139 6616 14280 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 14274 6604 14280 6616
rect 14332 6644 14338 6656
rect 14642 6644 14648 6656
rect 14332 6616 14648 6644
rect 14332 6604 14338 6616
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 15120 6644 15148 6684
rect 15810 6681 15822 6684
rect 15856 6712 15868 6715
rect 15930 6712 15936 6724
rect 15856 6684 15936 6712
rect 15856 6681 15868 6684
rect 15810 6675 15868 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16114 6672 16120 6724
rect 16172 6712 16178 6724
rect 17405 6715 17463 6721
rect 16172 6684 17080 6712
rect 16172 6672 16178 6684
rect 14792 6616 15148 6644
rect 14792 6604 14798 6616
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 17052 6653 17080 6684
rect 17405 6681 17417 6715
rect 17451 6712 17463 6715
rect 18322 6712 18328 6724
rect 17451 6684 18328 6712
rect 17451 6681 17463 6684
rect 17405 6675 17463 6681
rect 18322 6672 18328 6684
rect 18380 6672 18386 6724
rect 16945 6647 17003 6653
rect 16945 6644 16957 6647
rect 16264 6616 16957 6644
rect 16264 6604 16270 6616
rect 16945 6613 16957 6616
rect 16991 6613 17003 6647
rect 16945 6607 17003 6613
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18414 6644 18420 6656
rect 18095 6616 18420 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1762 6440 1768 6452
rect 1723 6412 1768 6440
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2464 6412 2789 6440
rect 2464 6400 2470 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 2777 6403 2835 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3660 6412 3985 6440
rect 3660 6400 3666 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 12250 6440 12256 6452
rect 3973 6403 4031 6409
rect 5000 6412 12256 6440
rect 2590 6332 2596 6384
rect 2648 6372 2654 6384
rect 4065 6375 4123 6381
rect 4065 6372 4077 6375
rect 2648 6344 4077 6372
rect 2648 6332 2654 6344
rect 4065 6341 4077 6344
rect 4111 6341 4123 6375
rect 4065 6335 4123 6341
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 5000 6372 5028 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12434 6440 12440 6452
rect 12395 6412 12440 6440
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13170 6440 13176 6452
rect 12820 6412 13176 6440
rect 12820 6372 12848 6412
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 14090 6440 14096 6452
rect 13495 6412 14096 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 15838 6440 15844 6452
rect 15580 6412 15844 6440
rect 4488 6344 4844 6372
rect 4488 6332 4494 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2222 6304 2228 6316
rect 2183 6276 2228 6304
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 4246 6304 4252 6316
rect 3191 6276 4252 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4816 6313 4844 6344
rect 4908 6344 5028 6372
rect 6012 6344 12848 6372
rect 14584 6375 14642 6381
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3602 6236 3608 6248
rect 3467 6208 3608 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4338 6236 4344 6248
rect 3927 6208 4344 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4908 6236 4936 6344
rect 5074 6313 5080 6316
rect 5068 6304 5080 6313
rect 4987 6276 5080 6304
rect 5068 6267 5080 6276
rect 5132 6304 5138 6316
rect 5350 6304 5356 6316
rect 5132 6276 5356 6304
rect 5074 6264 5080 6267
rect 5132 6264 5138 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5810 6264 5816 6316
rect 5868 6304 5874 6316
rect 6012 6304 6040 6344
rect 14584 6341 14596 6375
rect 14630 6372 14642 6375
rect 15580 6372 15608 6412
rect 15838 6400 15844 6412
rect 15896 6440 15902 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 15896 6412 16313 6440
rect 15896 6400 15902 6412
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 16301 6403 16359 6409
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6440 16911 6443
rect 18230 6440 18236 6452
rect 16899 6412 18236 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 18414 6440 18420 6452
rect 18375 6412 18420 6440
rect 18414 6400 18420 6412
rect 18472 6400 18478 6452
rect 14630 6344 15608 6372
rect 14630 6341 14642 6344
rect 14584 6335 14642 6341
rect 16390 6332 16396 6384
rect 16448 6372 16454 6384
rect 16448 6344 17448 6372
rect 16448 6332 16454 6344
rect 17420 6328 17448 6344
rect 5868 6276 6040 6304
rect 5868 6264 5874 6276
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6362 6304 6368 6316
rect 6236 6276 6368 6304
rect 6236 6264 6242 6276
rect 6362 6264 6368 6276
rect 6420 6304 6426 6316
rect 7357 6307 7415 6313
rect 7357 6304 7369 6307
rect 6420 6276 7369 6304
rect 6420 6264 6426 6276
rect 7357 6273 7369 6276
rect 7403 6273 7415 6307
rect 7357 6267 7415 6273
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9490 6313 9496 6316
rect 9484 6304 9496 6313
rect 8996 6276 9496 6304
rect 8996 6264 9002 6276
rect 9484 6267 9496 6276
rect 9490 6264 9496 6267
rect 9548 6264 9554 6316
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 10744 6276 11989 6304
rect 10744 6264 10750 6276
rect 11977 6273 11989 6276
rect 12023 6304 12035 6307
rect 12621 6307 12679 6313
rect 12023 6276 12434 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 4816 6208 4936 6236
rect 6457 6239 6515 6245
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6168 2743 6171
rect 3050 6168 3056 6180
rect 2731 6140 3056 6168
rect 2731 6137 2743 6140
rect 2685 6131 2743 6137
rect 3050 6128 3056 6140
rect 3108 6168 3114 6180
rect 4816 6168 4844 6208
rect 6457 6205 6469 6239
rect 6503 6236 6515 6239
rect 6638 6236 6644 6248
rect 6503 6208 6644 6236
rect 6503 6205 6515 6208
rect 6457 6199 6515 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6880 6208 7113 6236
rect 6880 6196 6886 6208
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 9214 6236 9220 6248
rect 9175 6208 9220 6236
rect 7101 6199 7159 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 11514 6236 11520 6248
rect 10284 6208 11520 6236
rect 10284 6196 10290 6208
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 12158 6236 12164 6248
rect 12119 6208 12164 6236
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 12406 6236 12434 6276
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12802 6304 12808 6316
rect 12667 6276 12808 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 12894 6264 12900 6316
rect 12952 6304 12958 6316
rect 13081 6308 13139 6313
rect 13004 6307 13139 6308
rect 13004 6304 13093 6307
rect 12952 6280 13093 6304
rect 12952 6276 13032 6280
rect 12952 6264 12958 6276
rect 13081 6273 13093 6280
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6304 14887 6307
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14875 6276 14933 6304
rect 14875 6273 14887 6276
rect 14829 6267 14887 6273
rect 14921 6273 14933 6276
rect 14967 6304 14979 6307
rect 15010 6304 15016 6316
rect 14967 6276 15016 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 12986 6236 12992 6248
rect 12406 6208 12992 6236
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 11333 6171 11391 6177
rect 3108 6140 4844 6168
rect 5736 6140 7052 6168
rect 3108 6128 3114 6140
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 2004 6072 2053 6100
rect 2004 6060 2010 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 2280 6072 2329 6100
rect 2280 6060 2286 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 2317 6063 2375 6069
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 3142 6100 3148 6112
rect 2648 6072 3148 6100
rect 2648 6060 2654 6072
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4430 6100 4436 6112
rect 4391 6072 4436 6100
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 4706 6100 4712 6112
rect 4663 6072 4712 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5166 6060 5172 6112
rect 5224 6100 5230 6112
rect 5736 6100 5764 6140
rect 6178 6100 6184 6112
rect 5224 6072 5764 6100
rect 6139 6072 6184 6100
rect 5224 6060 5230 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6546 6100 6552 6112
rect 6420 6072 6552 6100
rect 6420 6060 6426 6072
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6730 6100 6736 6112
rect 6691 6072 6736 6100
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 6914 6100 6920 6112
rect 6875 6072 6920 6100
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7024 6100 7052 6140
rect 8036 6140 8616 6168
rect 8036 6100 8064 6140
rect 7024 6072 8064 6100
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 8352 6072 8493 6100
rect 8352 6060 8358 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 8588 6100 8616 6140
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 11606 6168 11612 6180
rect 11379 6140 11612 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 13197 6168 13225 6267
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15188 6307 15246 6313
rect 15188 6273 15200 6307
rect 15234 6304 15246 6307
rect 16298 6304 16304 6316
rect 15234 6276 16304 6304
rect 15234 6273 15246 6276
rect 15188 6267 15246 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16531 6276 16681 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16669 6273 16681 6276
rect 16715 6304 16727 6307
rect 16850 6304 16856 6316
rect 16715 6276 16856 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 17420 6313 17724 6328
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 17092 6276 17233 6304
rect 17092 6264 17098 6276
rect 17221 6273 17233 6276
rect 17267 6273 17279 6307
rect 17420 6307 17739 6313
rect 17420 6300 17693 6307
rect 17221 6267 17279 6273
rect 17681 6273 17693 6300
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 17773 6308 17831 6313
rect 17773 6307 18000 6308
rect 17773 6273 17785 6307
rect 17819 6304 18000 6307
rect 18046 6304 18052 6316
rect 17819 6280 18052 6304
rect 17819 6273 17831 6280
rect 17972 6276 18052 6280
rect 17773 6267 17831 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 18230 6304 18236 6316
rect 18191 6276 18236 6304
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6205 17923 6239
rect 17865 6199 17923 6205
rect 12728 6140 13225 6168
rect 13357 6171 13415 6177
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 8588 6072 10609 6100
rect 8481 6063 8539 6069
rect 10597 6069 10609 6072
rect 10643 6100 10655 6103
rect 10686 6100 10692 6112
rect 10643 6072 10692 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11204 6072 11529 6100
rect 11204 6060 11210 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 11517 6063 11575 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 12728 6109 12756 6140
rect 13357 6137 13369 6171
rect 13403 6168 13415 6171
rect 13403 6140 13952 6168
rect 13403 6137 13415 6140
rect 13357 6131 13415 6137
rect 12713 6103 12771 6109
rect 12713 6100 12725 6103
rect 12676 6072 12725 6100
rect 12676 6060 12682 6072
rect 12713 6069 12725 6072
rect 12759 6069 12771 6103
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12713 6063 12771 6069
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13924 6100 13952 6140
rect 14090 6100 14096 6112
rect 13924 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 17034 6100 17040 6112
rect 16995 6072 17040 6100
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 17310 6100 17316 6112
rect 17271 6072 17316 6100
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 17880 6100 17908 6199
rect 17828 6072 17908 6100
rect 17828 6060 17834 6072
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 2866 5896 2872 5908
rect 2823 5868 2872 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 4246 5856 4252 5868
rect 4304 5896 4310 5908
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 4304 5868 5120 5896
rect 4304 5856 4310 5868
rect 3605 5831 3663 5837
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 4798 5828 4804 5840
rect 3651 5800 4804 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 2133 5763 2191 5769
rect 2133 5760 2145 5763
rect 1544 5732 2145 5760
rect 1544 5720 1550 5732
rect 2133 5729 2145 5732
rect 2179 5729 2191 5763
rect 2133 5723 2191 5729
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5760 2375 5763
rect 2682 5760 2688 5772
rect 2363 5732 2688 5760
rect 2363 5729 2375 5732
rect 2317 5723 2375 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3050 5760 3056 5772
rect 3011 5732 3056 5760
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 4522 5720 4528 5772
rect 4580 5720 4586 5772
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 4985 5763 5043 5769
rect 4985 5760 4997 5763
rect 4672 5732 4997 5760
rect 4672 5720 4678 5732
rect 4985 5729 4997 5732
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 3973 5711 4031 5717
rect 3973 5708 3985 5711
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 2409 5695 2467 5701
rect 2409 5692 2421 5695
rect 1995 5664 2421 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 2409 5661 2421 5664
rect 2455 5692 2467 5695
rect 3142 5692 3148 5704
rect 2455 5664 3148 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 3804 5692 3985 5708
rect 3476 5680 3985 5692
rect 3476 5664 3832 5680
rect 3973 5677 3985 5680
rect 4019 5677 4031 5711
rect 4540 5692 4568 5720
rect 4706 5692 4712 5704
rect 3973 5671 4031 5677
rect 4065 5671 4123 5677
rect 3476 5652 3482 5664
rect 4065 5637 4077 5671
rect 4111 5668 4123 5671
rect 4111 5640 4200 5668
rect 4540 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 5092 5692 5120 5868
rect 5184 5868 11989 5896
rect 5184 5769 5212 5868
rect 11977 5865 11989 5868
rect 12023 5896 12035 5899
rect 12342 5896 12348 5908
rect 12023 5868 12348 5896
rect 12023 5865 12035 5868
rect 11977 5859 12035 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 13320 5868 13553 5896
rect 13320 5856 13326 5868
rect 13541 5865 13553 5868
rect 13587 5896 13599 5899
rect 13587 5868 15424 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 5408 5800 6101 5828
rect 5408 5788 5414 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 12066 5828 12072 5840
rect 12027 5800 12072 5828
rect 6089 5791 6147 5797
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 15396 5828 15424 5868
rect 15470 5856 15476 5908
rect 15528 5896 15534 5908
rect 15565 5899 15623 5905
rect 15565 5896 15577 5899
rect 15528 5868 15577 5896
rect 15528 5856 15534 5868
rect 15565 5865 15577 5868
rect 15611 5865 15623 5899
rect 15565 5859 15623 5865
rect 16206 5856 16212 5908
rect 16264 5896 16270 5908
rect 16850 5896 16856 5908
rect 16264 5868 16856 5896
rect 16264 5856 16270 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 15930 5828 15936 5840
rect 15396 5800 15936 5828
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 16758 5788 16764 5840
rect 16816 5828 16822 5840
rect 17586 5828 17592 5840
rect 16816 5800 17592 5828
rect 16816 5788 16822 5800
rect 17586 5788 17592 5800
rect 17644 5828 17650 5840
rect 17644 5800 18368 5828
rect 17644 5788 17650 5800
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 5169 5723 5227 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 11606 5720 11612 5772
rect 11664 5760 11670 5772
rect 12250 5760 12256 5772
rect 11664 5732 12256 5760
rect 11664 5720 11670 5732
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 13449 5763 13507 5769
rect 13449 5729 13461 5763
rect 13495 5760 13507 5763
rect 13495 5732 14136 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5092 5664 5549 5692
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6822 5692 6828 5704
rect 6696 5664 6828 5692
rect 6696 5652 6702 5664
rect 6822 5652 6828 5664
rect 6880 5692 6886 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 6880 5664 7481 5692
rect 6880 5652 6886 5664
rect 7469 5661 7481 5664
rect 7515 5692 7527 5695
rect 8110 5692 8116 5704
rect 7515 5664 8116 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8168 5664 9137 5692
rect 8168 5652 8174 5664
rect 9125 5661 9137 5664
rect 9171 5692 9183 5695
rect 9214 5692 9220 5704
rect 9171 5664 9220 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9392 5695 9450 5701
rect 9392 5692 9404 5695
rect 9324 5664 9404 5692
rect 4111 5637 4123 5640
rect 1210 5584 1216 5636
rect 1268 5624 1274 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 1268 5596 3249 5624
rect 1268 5584 1274 5596
rect 3237 5593 3249 5596
rect 3283 5624 3295 5627
rect 3326 5624 3332 5636
rect 3283 5596 3332 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 4065 5631 4123 5637
rect 4172 5624 4200 5640
rect 4341 5627 4399 5633
rect 4341 5624 4353 5627
rect 3436 5596 3924 5624
rect 4172 5596 4353 5624
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 3436 5556 3464 5596
rect 3191 5528 3464 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3752 5528 3801 5556
rect 3752 5516 3758 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3896 5556 3924 5596
rect 4341 5593 4353 5596
rect 4387 5624 4399 5627
rect 4387 5596 5764 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 4356 5556 4384 5587
rect 3896 5528 4384 5556
rect 3789 5519 3847 5525
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 4488 5528 4537 5556
rect 4488 5516 4494 5528
rect 4525 5525 4537 5528
rect 4571 5525 4583 5559
rect 4525 5519 4583 5525
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 4893 5559 4951 5565
rect 4893 5556 4905 5559
rect 4672 5528 4905 5556
rect 4672 5516 4678 5528
rect 4893 5525 4905 5528
rect 4939 5525 4951 5559
rect 4893 5519 4951 5525
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5736 5565 5764 5596
rect 7098 5584 7104 5636
rect 7156 5624 7162 5636
rect 7202 5627 7260 5633
rect 7202 5624 7214 5627
rect 7156 5596 7214 5624
rect 7156 5584 7162 5596
rect 7202 5593 7214 5596
rect 7248 5593 7260 5627
rect 7202 5587 7260 5593
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 5040 5528 5365 5556
rect 5040 5516 5046 5528
rect 5353 5525 5365 5528
rect 5399 5525 5411 5559
rect 5353 5519 5411 5525
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 8202 5556 8208 5568
rect 5767 5528 8208 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 9232 5556 9260 5652
rect 9324 5636 9352 5664
rect 9392 5661 9404 5664
rect 9438 5692 9450 5695
rect 10226 5692 10232 5704
rect 9438 5664 10232 5692
rect 9438 5661 9450 5664
rect 9392 5655 9450 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 11330 5692 11336 5704
rect 10643 5664 11336 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 9306 5584 9312 5636
rect 9364 5584 9370 5636
rect 10612 5624 10640 5655
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 13906 5692 13912 5704
rect 13771 5664 13912 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 14108 5701 14136 5732
rect 16390 5720 16396 5772
rect 16448 5760 16454 5772
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 16448 5732 16681 5760
rect 16448 5720 16454 5732
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 18340 5769 18368 5800
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 17460 5732 17509 5760
rect 17460 5720 17466 5732
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14182 5692 14188 5704
rect 14139 5664 14188 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14182 5652 14188 5664
rect 14240 5692 14246 5704
rect 15102 5692 15108 5704
rect 14240 5664 15108 5692
rect 14240 5652 14246 5664
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 15304 5664 15761 5692
rect 9646 5596 10640 5624
rect 9646 5556 9674 5596
rect 10686 5584 10692 5636
rect 10744 5624 10750 5636
rect 10842 5627 10900 5633
rect 10842 5624 10854 5627
rect 10744 5596 10854 5624
rect 10744 5584 10750 5596
rect 10842 5593 10854 5596
rect 10888 5593 10900 5627
rect 13078 5624 13084 5636
rect 10842 5587 10900 5593
rect 12268 5596 13084 5624
rect 9232 5528 9674 5556
rect 10505 5559 10563 5565
rect 10505 5525 10517 5559
rect 10551 5556 10563 5559
rect 12268 5556 12296 5596
rect 13078 5584 13084 5596
rect 13136 5624 13142 5636
rect 13182 5627 13240 5633
rect 13182 5624 13194 5627
rect 13136 5596 13194 5624
rect 13136 5584 13142 5596
rect 13182 5593 13194 5596
rect 13228 5593 13240 5627
rect 13182 5587 13240 5593
rect 14360 5627 14418 5633
rect 14360 5593 14372 5627
rect 14406 5624 14418 5627
rect 15194 5624 15200 5636
rect 14406 5596 15200 5624
rect 14406 5593 14418 5596
rect 14360 5587 14418 5593
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 10551 5528 12296 5556
rect 10551 5525 10563 5528
rect 10505 5519 10563 5525
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 13722 5556 13728 5568
rect 12400 5528 13728 5556
rect 12400 5516 12406 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 15304 5556 15332 5664
rect 15749 5661 15761 5664
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 17310 5692 17316 5704
rect 16531 5664 17316 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 16577 5627 16635 5633
rect 15488 5596 16528 5624
rect 15488 5568 15516 5596
rect 15470 5556 15476 5568
rect 13955 5528 15332 5556
rect 15431 5528 15476 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 15838 5516 15844 5568
rect 15896 5556 15902 5568
rect 15933 5559 15991 5565
rect 15933 5556 15945 5559
rect 15896 5528 15945 5556
rect 15896 5516 15902 5528
rect 15933 5525 15945 5528
rect 15979 5525 15991 5559
rect 16114 5556 16120 5568
rect 16075 5528 16120 5556
rect 15933 5519 15991 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16500 5556 16528 5596
rect 16577 5593 16589 5627
rect 16623 5624 16635 5627
rect 17494 5624 17500 5636
rect 16623 5596 17500 5624
rect 16623 5593 16635 5596
rect 16577 5587 16635 5593
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 16758 5556 16764 5568
rect 16500 5528 16764 5556
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 16850 5516 16856 5568
rect 16908 5556 16914 5568
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 16908 5528 16957 5556
rect 16908 5516 16914 5528
rect 16945 5525 16957 5528
rect 16991 5525 17003 5559
rect 17310 5556 17316 5568
rect 17271 5528 17316 5556
rect 16945 5519 17003 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 17451 5528 17785 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 17773 5519 17831 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 18288 5528 18333 5556
rect 18288 5516 18294 5528
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3602 5352 3608 5364
rect 3191 5324 3608 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 3878 5312 3884 5364
rect 3936 5352 3942 5364
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3936 5324 3985 5352
rect 3936 5312 3942 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4111 5324 4445 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4798 5352 4804 5364
rect 4759 5324 4804 5352
rect 4433 5315 4491 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5352 4951 5355
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4939 5324 5273 5352
rect 4939 5321 4951 5324
rect 4893 5315 4951 5321
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 9306 5352 9312 5364
rect 8067 5324 9312 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 9493 5355 9551 5361
rect 9493 5352 9505 5355
rect 9456 5324 9505 5352
rect 9456 5312 9462 5324
rect 9493 5321 9505 5324
rect 9539 5321 9551 5355
rect 11974 5352 11980 5364
rect 9493 5315 9551 5321
rect 9646 5324 11980 5352
rect 1854 5244 1860 5296
rect 1912 5284 1918 5296
rect 3620 5284 3648 5312
rect 5629 5287 5687 5293
rect 5629 5284 5641 5287
rect 1912 5256 2360 5284
rect 3620 5256 5641 5284
rect 1912 5244 1918 5256
rect 1670 5216 1676 5228
rect 1631 5188 1676 5216
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2222 5216 2228 5228
rect 2087 5188 2228 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2332 5225 2360 5256
rect 5276 5228 5304 5256
rect 5629 5253 5641 5256
rect 5675 5253 5687 5287
rect 5629 5247 5687 5253
rect 6270 5244 6276 5296
rect 6328 5284 6334 5296
rect 6886 5287 6944 5293
rect 6886 5284 6898 5287
rect 6328 5256 6898 5284
rect 6328 5244 6334 5256
rect 6886 5253 6898 5256
rect 6932 5253 6944 5287
rect 6886 5247 6944 5253
rect 7374 5244 7380 5296
rect 7432 5284 7438 5296
rect 9646 5284 9674 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16298 5352 16304 5364
rect 15887 5324 16304 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 17368 5324 17417 5352
rect 17368 5312 17374 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 18230 5352 18236 5364
rect 18191 5324 18236 5352
rect 17405 5315 17463 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18380 5324 18425 5352
rect 18380 5312 18386 5324
rect 11330 5284 11336 5296
rect 7432 5256 9674 5284
rect 9968 5256 11336 5284
rect 7432 5244 7438 5256
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2590 5216 2596 5228
rect 2551 5188 2596 5216
rect 2317 5179 2375 5185
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 5258 5176 5264 5228
rect 5316 5176 5322 5228
rect 6638 5216 6644 5228
rect 6599 5188 6644 5216
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 8110 5216 8116 5228
rect 7248 5188 7972 5216
rect 8071 5188 8116 5216
rect 7248 5176 7254 5188
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3237 5151 3295 5157
rect 3237 5148 3249 5151
rect 2924 5120 3249 5148
rect 2924 5108 2930 5120
rect 3237 5117 3249 5120
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 3878 5148 3884 5160
rect 3375 5120 3884 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4890 5148 4896 5160
rect 4295 5120 4896 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5074 5148 5080 5160
rect 5035 5120 5080 5148
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5718 5148 5724 5160
rect 5679 5120 5724 5148
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5117 5871 5151
rect 7944 5148 7972 5188
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 9968 5225 9996 5256
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 14182 5284 14188 5296
rect 12912 5256 14188 5284
rect 10226 5225 10232 5228
rect 8369 5219 8427 5225
rect 8369 5216 8381 5219
rect 8220 5188 8381 5216
rect 8220 5148 8248 5188
rect 8369 5185 8381 5188
rect 8415 5185 8427 5219
rect 8369 5179 8427 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 10220 5216 10232 5225
rect 10187 5188 10232 5216
rect 9953 5179 10011 5185
rect 10220 5179 10232 5188
rect 10226 5176 10232 5179
rect 10284 5176 10290 5228
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 12912 5225 12940 5256
rect 14182 5244 14188 5256
rect 14240 5284 14246 5296
rect 14240 5256 14412 5284
rect 14240 5244 14246 5256
rect 12630 5219 12688 5225
rect 12630 5216 12642 5219
rect 10744 5188 12642 5216
rect 10744 5176 10750 5188
rect 12630 5185 12642 5188
rect 12676 5185 12688 5219
rect 12630 5179 12688 5185
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 14384 5225 14412 5256
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17494 5284 17500 5296
rect 17000 5256 17500 5284
rect 17000 5244 17006 5256
rect 17494 5244 17500 5256
rect 17552 5284 17558 5296
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 17552 5256 17785 5284
rect 17552 5244 17558 5256
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 14102 5219 14160 5225
rect 14102 5216 14114 5219
rect 13780 5188 14114 5216
rect 13780 5176 13786 5188
rect 14102 5185 14114 5188
rect 14148 5185 14160 5219
rect 14102 5179 14160 5185
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14415 5188 14473 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14728 5219 14786 5225
rect 14728 5185 14740 5219
rect 14774 5216 14786 5219
rect 15654 5216 15660 5228
rect 14774 5188 15660 5216
rect 14774 5185 14786 5188
rect 14728 5179 14786 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 7944 5120 8248 5148
rect 5813 5111 5871 5117
rect 2038 5040 2044 5092
rect 2096 5080 2102 5092
rect 2409 5083 2467 5089
rect 2409 5080 2421 5083
rect 2096 5052 2421 5080
rect 2096 5040 2102 5052
rect 2409 5049 2421 5052
rect 2455 5049 2467 5083
rect 2409 5043 2467 5049
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 2958 5080 2964 5092
rect 2648 5052 2964 5080
rect 2648 5040 2654 5052
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 3476 5052 3832 5080
rect 3476 5040 3482 5052
rect 1486 4972 1492 5024
rect 1544 5012 1550 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1544 4984 1869 5012
rect 1544 4972 1550 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 2222 5012 2228 5024
rect 2179 4984 2228 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 3605 5015 3663 5021
rect 2832 4984 2877 5012
rect 2832 4972 2838 4984
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 3694 5012 3700 5024
rect 3651 4984 3700 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 3804 5012 3832 5052
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4614 5080 4620 5092
rect 4212 5052 4620 5080
rect 4212 5040 4218 5052
rect 4614 5040 4620 5052
rect 4672 5080 4678 5092
rect 5442 5080 5448 5092
rect 4672 5052 5448 5080
rect 4672 5040 4678 5052
rect 5442 5040 5448 5052
rect 5500 5080 5506 5092
rect 5828 5080 5856 5111
rect 5500 5052 5856 5080
rect 6181 5083 6239 5089
rect 5500 5040 5506 5052
rect 6181 5049 6193 5083
rect 6227 5080 6239 5083
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 6227 5052 6684 5080
rect 6227 5049 6239 5052
rect 6181 5043 6239 5049
rect 6196 5012 6224 5043
rect 3804 4984 6224 5012
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 6328 4984 6377 5012
rect 6328 4972 6334 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6656 5012 6684 5052
rect 10888 5052 11529 5080
rect 8754 5012 8760 5024
rect 6656 4984 8760 5012
rect 6365 4975 6423 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10888 5012 10916 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 16117 5083 16175 5089
rect 16117 5049 16129 5083
rect 16163 5080 16175 5083
rect 16500 5080 16528 5179
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16632 5188 17049 5216
rect 16632 5176 16638 5188
rect 17037 5185 17049 5188
rect 17083 5216 17095 5219
rect 17865 5219 17923 5225
rect 17083 5188 17724 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 16758 5148 16764 5160
rect 16719 5120 16764 5148
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16942 5148 16948 5160
rect 16903 5120 16948 5148
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 17589 5151 17647 5157
rect 17589 5148 17601 5151
rect 17368 5120 17601 5148
rect 17368 5108 17374 5120
rect 17589 5117 17601 5120
rect 17635 5117 17647 5151
rect 17696 5148 17724 5188
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 18598 5216 18604 5228
rect 17911 5188 18604 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 18966 5148 18972 5160
rect 17696 5120 18972 5148
rect 17589 5111 17647 5117
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 18322 5080 18328 5092
rect 16163 5052 16436 5080
rect 16500 5052 18328 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 9640 4984 10916 5012
rect 11333 5015 11391 5021
rect 9640 4972 9646 4984
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 11422 5012 11428 5024
rect 11379 4984 11428 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12989 5015 13047 5021
rect 12989 5012 13001 5015
rect 12032 4984 13001 5012
rect 12032 4972 12038 4984
rect 12989 4981 13001 4984
rect 13035 4981 13047 5015
rect 16298 5012 16304 5024
rect 16259 4984 16304 5012
rect 12989 4975 13047 4981
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 16408 5012 16436 5052
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 18230 5012 18236 5024
rect 16408 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 2866 4808 2872 4820
rect 2827 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 4522 4808 4528 4820
rect 3936 4780 4528 4808
rect 3936 4768 3942 4780
rect 4522 4768 4528 4780
rect 4580 4808 4586 4820
rect 4798 4808 4804 4820
rect 4580 4780 4804 4808
rect 4580 4768 4586 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6086 4808 6092 4820
rect 5859 4780 6092 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 6880 4780 7236 4808
rect 6880 4768 6886 4780
rect 1765 4743 1823 4749
rect 1765 4709 1777 4743
rect 1811 4709 1823 4743
rect 3418 4740 3424 4752
rect 3331 4712 3424 4740
rect 1765 4703 1823 4709
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 1780 4604 1808 4703
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 2774 4672 2780 4684
rect 2363 4644 2780 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 1946 4604 1952 4616
rect 1719 4576 1808 4604
rect 1907 4576 1952 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2240 4604 2268 4635
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3344 4681 3372 4712
rect 3418 4700 3424 4712
rect 3476 4740 3482 4752
rect 4062 4740 4068 4752
rect 3476 4712 4068 4740
rect 3476 4700 3482 4712
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 7208 4681 7236 4780
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8076 4780 9045 4808
rect 8076 4768 8082 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 14734 4808 14740 4820
rect 11480 4780 14740 4808
rect 11480 4768 11486 4780
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15252 4780 15516 4808
rect 15252 4768 15258 4780
rect 13722 4700 13728 4752
rect 13780 4740 13786 4752
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 13780 4712 14105 4740
rect 13780 4700 13786 4712
rect 14093 4709 14105 4712
rect 14139 4709 14151 4743
rect 14093 4703 14151 4709
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 7193 4675 7251 4681
rect 3559 4644 4752 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 2590 4604 2596 4616
rect 2240 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3050 4564 3056 4616
rect 3108 4604 3114 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3108 4576 3249 4604
rect 3108 4564 3114 4576
rect 3237 4573 3249 4576
rect 3283 4604 3295 4607
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3283 4576 3985 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 4212 4576 4261 4604
rect 4212 4564 4218 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4724 4604 4752 4644
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 7239 4644 7389 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4672 10471 4675
rect 11330 4672 11336 4684
rect 10459 4644 11336 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 11330 4632 11336 4644
rect 11388 4672 11394 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11388 4644 11713 4672
rect 11388 4632 11394 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 5074 4604 5080 4616
rect 4724 4576 5080 4604
rect 4249 4567 4307 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5442 4564 5448 4616
rect 5500 4613 5506 4616
rect 5500 4604 5512 4613
rect 5721 4607 5779 4613
rect 5500 4576 5545 4604
rect 5500 4567 5512 4576
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6638 4604 6644 4616
rect 5767 4576 6644 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 5500 4564 5506 4567
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 6926 4607 6984 4613
rect 6926 4573 6938 4607
rect 6972 4604 6984 4607
rect 6972 4576 7052 4604
rect 6972 4573 6984 4576
rect 6926 4567 6984 4573
rect 7024 4548 7052 4576
rect 10134 4564 10140 4616
rect 10192 4613 10198 4616
rect 10192 4604 10204 4613
rect 10594 4604 10600 4616
rect 10192 4576 10456 4604
rect 10555 4576 10600 4604
rect 10192 4567 10204 4576
rect 10192 4564 10198 4567
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 6362 4536 6368 4548
rect 3200 4508 6368 4536
rect 3200 4496 3206 4508
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 7006 4496 7012 4548
rect 7064 4496 7070 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 7622 4539 7680 4545
rect 7622 4536 7634 4539
rect 7340 4508 7634 4536
rect 7340 4496 7346 4508
rect 7622 4505 7634 4508
rect 7668 4505 7680 4539
rect 9582 4536 9588 4548
rect 7622 4499 7680 4505
rect 8772 4508 9588 4536
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 2406 4468 2412 4480
rect 2367 4440 2412 4468
rect 2406 4428 2412 4440
rect 2464 4428 2470 4480
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3789 4471 3847 4477
rect 2832 4440 2877 4468
rect 2832 4428 2838 4440
rect 3789 4437 3801 4471
rect 3835 4468 3847 4471
rect 3878 4468 3884 4480
rect 3835 4440 3884 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4062 4468 4068 4480
rect 4023 4440 4068 4468
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4341 4471 4399 4477
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 4706 4468 4712 4480
rect 4387 4440 4712 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4706 4428 4712 4440
rect 4764 4468 4770 4480
rect 5166 4468 5172 4480
rect 4764 4440 5172 4468
rect 4764 4428 4770 4440
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 7024 4468 7052 4496
rect 7466 4468 7472 4480
rect 7024 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 8772 4477 8800 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 10428 4536 10456 4576
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 11848 4576 13277 4604
rect 11848 4564 11854 4576
rect 13265 4573 13277 4576
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 13633 4607 13691 4613
rect 13633 4573 13645 4607
rect 13679 4573 13691 4607
rect 14108 4604 14136 4703
rect 15488 4681 15516 4780
rect 16758 4768 16764 4820
rect 16816 4808 16822 4820
rect 17034 4808 17040 4820
rect 16816 4780 17040 4808
rect 16816 4768 16822 4780
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 17957 4811 18015 4817
rect 17957 4777 17969 4811
rect 18003 4808 18015 4811
rect 18138 4808 18144 4820
rect 18003 4780 18144 4808
rect 18003 4777 18015 4780
rect 17957 4771 18015 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18414 4808 18420 4820
rect 18375 4780 18420 4808
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 16390 4740 16396 4752
rect 15620 4712 16396 4740
rect 15620 4700 15626 4712
rect 16390 4700 16396 4712
rect 16448 4740 16454 4752
rect 16448 4712 16988 4740
rect 16448 4700 16454 4712
rect 15473 4675 15531 4681
rect 15473 4641 15485 4675
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 15657 4675 15715 4681
rect 15657 4641 15669 4675
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4672 15899 4675
rect 16850 4672 16856 4684
rect 15887 4644 16856 4672
rect 15887 4641 15899 4644
rect 15841 4635 15899 4641
rect 15672 4604 15700 4635
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 16960 4681 16988 4712
rect 16945 4675 17003 4681
rect 16945 4641 16957 4675
rect 16991 4641 17003 4675
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 16945 4635 17003 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4672 17555 4675
rect 17862 4672 17868 4684
rect 17543 4644 17868 4672
rect 17543 4641 17555 4644
rect 17497 4635 17555 4641
rect 14108 4576 15700 4604
rect 13633 4567 13691 4573
rect 11514 4536 11520 4548
rect 10428 4508 11520 4536
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 11968 4539 12026 4545
rect 11968 4505 11980 4539
rect 12014 4536 12026 4539
rect 12014 4508 12204 4536
rect 12014 4505 12026 4508
rect 11968 4499 12026 4505
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4437 8815 4471
rect 12176 4468 12204 4508
rect 12250 4496 12256 4548
rect 12308 4536 12314 4548
rect 13648 4536 13676 4567
rect 15746 4564 15752 4616
rect 15804 4604 15810 4616
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15804 4576 15945 4604
rect 15804 4564 15810 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 17512 4604 17540 4635
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4672 18199 4675
rect 19058 4672 19064 4684
rect 18187 4644 19064 4672
rect 18187 4641 18199 4644
rect 18141 4635 18199 4641
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 17184 4576 17540 4604
rect 17589 4607 17647 4613
rect 17184 4564 17190 4576
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 17678 4604 17684 4616
rect 17635 4576 17684 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 18104 4576 18245 4604
rect 18104 4564 18110 4576
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 15102 4536 15108 4548
rect 12308 4508 13676 4536
rect 13740 4508 15108 4536
rect 12308 4496 12314 4508
rect 12434 4468 12440 4480
rect 12176 4440 12440 4468
rect 8757 4431 8815 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 13078 4468 13084 4480
rect 13039 4440 13084 4468
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13740 4468 13768 4508
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 15228 4539 15286 4545
rect 15228 4505 15240 4539
rect 15274 4536 15286 4539
rect 16022 4536 16028 4548
rect 15274 4508 16028 4536
rect 15274 4505 15286 4508
rect 15228 4499 15286 4505
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 16761 4539 16819 4545
rect 16761 4505 16773 4539
rect 16807 4536 16819 4539
rect 17402 4536 17408 4548
rect 16807 4508 17408 4536
rect 16807 4505 16819 4508
rect 16761 4499 16819 4505
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 13495 4440 13768 4468
rect 13817 4471 13875 4477
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13817 4437 13829 4471
rect 13863 4468 13875 4471
rect 15930 4468 15936 4480
rect 13863 4440 15936 4468
rect 13863 4437 13875 4440
rect 13817 4431 13875 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 16390 4428 16396 4480
rect 16448 4468 16454 4480
rect 16448 4440 16493 4468
rect 16448 4428 16454 4440
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 16908 4440 16953 4468
rect 16908 4428 16914 4440
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 1302 4224 1308 4276
rect 1360 4264 1366 4276
rect 2590 4264 2596 4276
rect 1360 4236 2596 4264
rect 1360 4224 1366 4236
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3513 4267 3571 4273
rect 3513 4264 3525 4267
rect 3108 4236 3525 4264
rect 3108 4224 3114 4236
rect 3513 4233 3525 4236
rect 3559 4264 3571 4267
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 3559 4236 4353 4264
rect 3559 4233 3571 4236
rect 3513 4227 3571 4233
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 4709 4267 4767 4273
rect 4709 4233 4721 4267
rect 4755 4264 4767 4267
rect 5718 4264 5724 4276
rect 4755 4236 5724 4264
rect 4755 4233 4767 4236
rect 4709 4227 4767 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 6181 4267 6239 4273
rect 6181 4233 6193 4267
rect 6227 4264 6239 4267
rect 11790 4264 11796 4276
rect 6227 4236 9674 4264
rect 11751 4236 11796 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 3418 4196 3424 4208
rect 2240 4168 2452 4196
rect 3379 4168 3424 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1854 4128 1860 4140
rect 1719 4100 1860 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2240 4060 2268 4168
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2424 4128 2452 4168
rect 3418 4156 3424 4168
rect 3476 4196 3482 4208
rect 4249 4199 4307 4205
rect 4249 4196 4261 4199
rect 3476 4168 4261 4196
rect 3476 4156 3482 4168
rect 4249 4165 4261 4168
rect 4295 4165 4307 4199
rect 4249 4159 4307 4165
rect 4522 4156 4528 4208
rect 4580 4196 4586 4208
rect 6196 4196 6224 4227
rect 4580 4168 6224 4196
rect 4580 4156 4586 4168
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 8076 4168 8524 4196
rect 8076 4156 8082 4168
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2424 4100 2605 4128
rect 2317 4091 2375 4097
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 2593 4091 2651 4097
rect 2056 4032 2268 4060
rect 2056 4004 2084 4032
rect 1486 3992 1492 4004
rect 1447 3964 1492 3992
rect 1486 3952 1492 3964
rect 1544 3952 1550 4004
rect 2038 3952 2044 4004
rect 2096 3952 2102 4004
rect 2332 3992 2360 4091
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 4706 4128 4712 4140
rect 4172 4100 4712 4128
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 4172 4069 4200 4100
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 5074 4137 5080 4140
rect 5068 4128 5080 4137
rect 5035 4100 5080 4128
rect 5068 4091 5080 4100
rect 5074 4088 5080 4091
rect 5132 4088 5138 4140
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5960 4100 6377 4128
rect 5960 4088 5966 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 7857 4131 7915 4137
rect 7857 4128 7869 4131
rect 6604 4100 7869 4128
rect 6604 4088 6610 4100
rect 7857 4097 7869 4100
rect 7903 4128 7915 4131
rect 8113 4131 8171 4137
rect 7903 4100 8064 4128
rect 7903 4097 7915 4100
rect 7857 4091 7915 4097
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 2556 4032 2789 4060
rect 2556 4020 2562 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2777 4023 2835 4029
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 8036 4060 8064 4100
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8202 4128 8208 4140
rect 8159 4100 8208 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8496 4128 8524 4168
rect 9502 4131 9560 4137
rect 9502 4128 9514 4131
rect 8496 4100 9514 4128
rect 9502 4097 9514 4100
rect 9548 4097 9560 4131
rect 9646 4128 9674 4236
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12069 4267 12127 4273
rect 12069 4233 12081 4267
rect 12115 4264 12127 4267
rect 12250 4264 12256 4276
rect 12115 4236 12256 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 15562 4264 15568 4276
rect 13136 4236 15568 4264
rect 13136 4224 13142 4236
rect 15562 4224 15568 4236
rect 15620 4224 15626 4276
rect 15841 4267 15899 4273
rect 15841 4233 15853 4267
rect 15887 4264 15899 4267
rect 16390 4264 16396 4276
rect 15887 4236 16396 4264
rect 15887 4233 15899 4236
rect 15841 4227 15899 4233
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17129 4267 17187 4273
rect 17129 4264 17141 4267
rect 17000 4236 17141 4264
rect 17000 4224 17006 4236
rect 17129 4233 17141 4236
rect 17175 4233 17187 4267
rect 17129 4227 17187 4233
rect 18417 4267 18475 4273
rect 18417 4233 18429 4267
rect 18463 4264 18475 4267
rect 18506 4264 18512 4276
rect 18463 4236 18512 4264
rect 18463 4233 18475 4236
rect 18417 4227 18475 4233
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 11330 4196 11336 4208
rect 9876 4168 11336 4196
rect 9876 4137 9904 4168
rect 11330 4156 11336 4168
rect 11388 4196 11394 4208
rect 15194 4196 15200 4208
rect 11388 4168 13584 4196
rect 11388 4156 11394 4168
rect 9769 4131 9827 4137
rect 9646 4100 9720 4128
rect 9502 4091 9560 4097
rect 8404 4060 8432 4088
rect 8036 4032 8432 4060
rect 9692 4060 9720 4100
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9815 4100 9873 4128
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 10117 4131 10175 4137
rect 10117 4128 10129 4131
rect 9861 4091 9919 4097
rect 9968 4100 10129 4128
rect 9968 4060 9996 4100
rect 10117 4097 10129 4100
rect 10163 4097 10175 4131
rect 10117 4091 10175 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11422 4128 11428 4140
rect 11296 4100 11428 4128
rect 11296 4088 11302 4100
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4128 11667 4131
rect 11698 4128 11704 4140
rect 11655 4100 11704 4128
rect 11655 4097 11667 4100
rect 11609 4091 11667 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12452 4137 12480 4168
rect 13556 4140 13584 4168
rect 14108 4168 15200 4196
rect 12710 4137 12716 4140
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 12483 4100 12517 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 12704 4091 12716 4137
rect 12768 4128 12774 4140
rect 12768 4100 12804 4128
rect 9692 4032 9996 4060
rect 4801 4023 4859 4029
rect 3142 3992 3148 4004
rect 2332 3964 3148 3992
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3344 3992 3372 4023
rect 4706 3992 4712 4004
rect 3344 3964 4712 3992
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 2004 3896 2145 3924
rect 2004 3884 2010 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2372 3896 2421 3924
rect 2372 3884 2378 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 3881 3927 3939 3933
rect 2924 3896 2969 3924
rect 2924 3884 2930 3896
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4246 3924 4252 3936
rect 3927 3896 4252 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4816 3924 4844 4023
rect 6733 3995 6791 4001
rect 6733 3961 6745 3995
rect 6779 3992 6791 3995
rect 7006 3992 7012 4004
rect 6779 3964 7012 3992
rect 6779 3961 6791 3964
rect 6733 3955 6791 3961
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 8168 3964 8401 3992
rect 8168 3952 8174 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 11606 3992 11612 4004
rect 8389 3955 8447 3961
rect 10796 3964 11612 3992
rect 5718 3924 5724 3936
rect 4816 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6328 3896 6561 3924
rect 6328 3884 6334 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 8297 3927 8355 3933
rect 8297 3893 8309 3927
rect 8343 3924 8355 3927
rect 8754 3924 8760 3936
rect 8343 3896 8760 3924
rect 8343 3893 8355 3896
rect 8297 3887 8355 3893
rect 8754 3884 8760 3896
rect 8812 3924 8818 3936
rect 10796 3924 10824 3964
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 12176 3992 12204 4091
rect 12710 4088 12716 4091
rect 12768 4088 12774 4100
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 14108 4137 14136 4168
rect 15194 4156 15200 4168
rect 15252 4156 15258 4208
rect 15933 4199 15991 4205
rect 15933 4165 15945 4199
rect 15979 4196 15991 4199
rect 16114 4196 16120 4208
rect 15979 4168 16120 4196
rect 15979 4165 15991 4168
rect 15933 4159 15991 4165
rect 16114 4156 16120 4168
rect 16172 4156 16178 4208
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 16816 4168 17540 4196
rect 16816 4156 16822 4168
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13596 4100 14105 4128
rect 13596 4088 13602 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14349 4131 14407 4137
rect 14349 4128 14361 4131
rect 14093 4091 14151 4097
rect 14200 4100 14361 4128
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14200 4060 14228 4100
rect 14349 4097 14361 4100
rect 14395 4097 14407 4131
rect 14349 4091 14407 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17218 4128 17224 4140
rect 17083 4100 17224 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17512 4137 17540 4168
rect 17586 4156 17592 4208
rect 17644 4196 17650 4208
rect 17644 4168 17689 4196
rect 17644 4156 17650 4168
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4097 18199 4131
rect 18141 4091 18199 4097
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18690 4128 18696 4140
rect 18279 4100 18696 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 13872 4032 14228 4060
rect 13872 4020 13878 4032
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 15654 4060 15660 4072
rect 15344 4032 15516 4060
rect 15615 4032 15660 4060
rect 15344 4020 15350 4032
rect 15488 4001 15516 4032
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 16264 4032 16405 4060
rect 16264 4020 16270 4032
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 17310 4060 17316 4072
rect 16393 4023 16451 4029
rect 16776 4032 17316 4060
rect 15473 3995 15531 4001
rect 12176 3964 12480 3992
rect 11238 3924 11244 3936
rect 8812 3896 10824 3924
rect 11199 3896 11244 3924
rect 8812 3884 8818 3896
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 12342 3924 12348 3936
rect 12303 3896 12348 3924
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12452 3924 12480 3964
rect 13372 3964 14044 3992
rect 13372 3924 13400 3964
rect 13814 3924 13820 3936
rect 12452 3896 13400 3924
rect 13775 3896 13820 3924
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14016 3933 14044 3964
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 16776 3992 16804 4032
rect 17310 4020 17316 4032
rect 17368 4060 17374 4072
rect 17681 4063 17739 4069
rect 17681 4060 17693 4063
rect 17368 4032 17693 4060
rect 17368 4020 17374 4032
rect 17681 4029 17693 4032
rect 17727 4029 17739 4063
rect 18156 4060 18184 4091
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18874 4060 18880 4072
rect 18156 4032 18880 4060
rect 17681 4023 17739 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 15519 3964 16804 3992
rect 16853 3995 16911 4001
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 17034 3992 17040 4004
rect 16899 3964 17040 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 17034 3952 17040 3964
rect 17092 3952 17098 4004
rect 17954 3992 17960 4004
rect 17915 3964 17960 3992
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 15286 3924 15292 3936
rect 14047 3896 15292 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 4154 3720 4160 3732
rect 3651 3692 4160 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4706 3680 4712 3732
rect 4764 3720 4770 3732
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 4764 3692 6653 3720
rect 4764 3680 4770 3692
rect 6641 3689 6653 3692
rect 6687 3720 6699 3723
rect 8570 3720 8576 3732
rect 6687 3692 8576 3720
rect 6687 3689 6699 3692
rect 6641 3683 6699 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 11054 3720 11060 3732
rect 8772 3692 11060 3720
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3652 2835 3655
rect 6546 3652 6552 3664
rect 2823 3624 4844 3652
rect 6507 3624 6552 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 1946 3584 1952 3596
rect 1688 3556 1952 3584
rect 1688 3525 1716 3556
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 3050 3584 3056 3596
rect 3011 3556 3056 3584
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 4430 3584 4436 3596
rect 3384 3556 4436 3584
rect 3384 3544 3390 3556
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 4522 3544 4528 3596
rect 4580 3584 4586 3596
rect 4580 3556 4625 3584
rect 4580 3544 4586 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2133 3519 2191 3525
rect 1820 3488 1865 3516
rect 1820 3476 1826 3488
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2222 3516 2228 3528
rect 2179 3488 2228 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2682 3516 2688 3528
rect 2639 3488 2688 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3145 3519 3203 3525
rect 3145 3516 3157 3519
rect 2832 3488 3157 3516
rect 2832 3476 2838 3488
rect 3145 3485 3157 3488
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3510 3516 3516 3528
rect 3283 3488 3516 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 3927 3488 4292 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4264 3448 4292 3488
rect 4338 3476 4344 3528
rect 4396 3516 4402 3528
rect 4816 3525 4844 3624
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8202 3584 8208 3596
rect 8067 3556 8208 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8404 3556 8616 3584
rect 4801 3519 4859 3525
rect 4396 3488 4476 3516
rect 4396 3476 4402 3488
rect 4448 3457 4476 3488
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5718 3516 5724 3528
rect 5215 3488 5724 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5718 3476 5724 3488
rect 5776 3516 5782 3528
rect 6178 3516 6184 3528
rect 5776 3488 6184 3516
rect 5776 3476 5782 3488
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 8404 3525 8432 3556
rect 7765 3519 7823 3525
rect 7765 3485 7777 3519
rect 7811 3516 7823 3519
rect 8382 3519 8440 3525
rect 7811 3488 8248 3516
rect 7811 3485 7823 3488
rect 7765 3479 7823 3485
rect 4433 3451 4491 3457
rect 2746 3420 4016 3448
rect 4264 3420 4384 3448
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 2280 3352 2329 3380
rect 2280 3340 2286 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 2406 3340 2412 3392
rect 2464 3380 2470 3392
rect 2746 3380 2774 3420
rect 3988 3389 4016 3420
rect 4356 3392 4384 3420
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4706 3448 4712 3460
rect 4479 3420 4712 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 4890 3408 4896 3460
rect 4948 3448 4954 3460
rect 5414 3451 5472 3457
rect 5414 3448 5426 3451
rect 4948 3420 5426 3448
rect 4948 3408 4954 3420
rect 5414 3417 5426 3420
rect 5460 3448 5472 3451
rect 8110 3448 8116 3460
rect 5460 3420 8116 3448
rect 5460 3417 5472 3420
rect 5414 3411 5472 3417
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8220 3448 8248 3488
rect 8382 3485 8394 3519
rect 8428 3485 8440 3519
rect 8382 3479 8440 3485
rect 8478 3476 8484 3528
rect 8536 3476 8542 3528
rect 8496 3448 8524 3476
rect 8220 3420 8524 3448
rect 8588 3448 8616 3556
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 8772 3516 8800 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 11440 3692 12173 3720
rect 9953 3655 10011 3661
rect 9953 3621 9965 3655
rect 9999 3652 10011 3655
rect 10318 3652 10324 3664
rect 9999 3624 10324 3652
rect 9999 3621 10011 3624
rect 9953 3615 10011 3621
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 11330 3584 11336 3596
rect 11291 3556 11336 3584
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 9122 3516 9128 3528
rect 8711 3488 8800 3516
rect 9083 3488 9128 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9398 3516 9404 3528
rect 9359 3488 9404 3516
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 9766 3516 9772 3528
rect 9631 3488 9772 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 11440 3516 11468 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 12161 3683 12219 3689
rect 15194 3680 15200 3732
rect 15252 3720 15258 3732
rect 15252 3692 15516 3720
rect 15252 3680 15258 3692
rect 11701 3655 11759 3661
rect 11701 3621 11713 3655
rect 11747 3652 11759 3655
rect 12342 3652 12348 3664
rect 11747 3624 12348 3652
rect 11747 3621 11759 3624
rect 11701 3615 11759 3621
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12526 3584 12532 3596
rect 11532 3556 12532 3584
rect 11532 3525 11560 3556
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 13538 3584 13544 3596
rect 13499 3556 13544 3584
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 15488 3593 15516 3692
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 16945 3723 17003 3729
rect 16945 3720 16957 3723
rect 15804 3692 16957 3720
rect 15804 3680 15810 3692
rect 16945 3689 16957 3692
rect 16991 3689 17003 3723
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 16945 3683 17003 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 17460 3692 17509 3720
rect 17460 3680 17466 3692
rect 17497 3689 17509 3692
rect 17543 3689 17555 3723
rect 18322 3720 18328 3732
rect 18283 3692 18328 3720
rect 17497 3683 17555 3689
rect 18322 3680 18328 3692
rect 18380 3680 18386 3732
rect 17770 3612 17776 3664
rect 17828 3652 17834 3664
rect 17828 3624 18092 3652
rect 17828 3612 17834 3624
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 15565 3587 15623 3593
rect 15565 3584 15577 3587
rect 15519 3556 15577 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 15565 3553 15577 3556
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 18064 3593 18092 3624
rect 17957 3587 18015 3593
rect 17957 3584 17969 3587
rect 17736 3556 17969 3584
rect 17736 3544 17742 3556
rect 17957 3553 17969 3556
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3553 18107 3587
rect 18782 3584 18788 3596
rect 18049 3547 18107 3553
rect 18156 3556 18788 3584
rect 9876 3488 11468 3516
rect 11517 3519 11575 3525
rect 8588 3420 9260 3448
rect 2464 3352 2774 3380
rect 3973 3383 4031 3389
rect 2464 3340 2470 3352
rect 3973 3349 3985 3383
rect 4019 3349 4031 3383
rect 4338 3380 4344 3392
rect 4299 3352 4344 3380
rect 3973 3343 4031 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 4985 3383 5043 3389
rect 4985 3380 4997 3383
rect 4580 3352 4997 3380
rect 4580 3340 4586 3352
rect 4985 3349 4997 3352
rect 5031 3349 5043 3383
rect 4985 3343 5043 3349
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 7926 3380 7932 3392
rect 5224 3352 7932 3380
rect 5224 3340 5230 3352
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 8076 3352 8217 3380
rect 8076 3340 8082 3352
rect 8205 3349 8217 3352
rect 8251 3349 8263 3383
rect 8205 3343 8263 3349
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8481 3383 8539 3389
rect 8481 3380 8493 3383
rect 8444 3352 8493 3380
rect 8444 3340 8450 3352
rect 8481 3349 8493 3352
rect 8527 3349 8539 3383
rect 8481 3343 8539 3349
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9232 3389 9260 3420
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 9876 3448 9904 3488
rect 11517 3485 11529 3519
rect 11563 3485 11575 3519
rect 11974 3516 11980 3528
rect 11517 3479 11575 3485
rect 11808 3488 11980 3516
rect 9364 3420 9904 3448
rect 11088 3451 11146 3457
rect 9364 3408 9370 3420
rect 11088 3417 11100 3451
rect 11134 3448 11146 3451
rect 11808 3448 11836 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3516 12127 3519
rect 12894 3516 12900 3528
rect 12115 3488 12900 3516
rect 12115 3485 12127 3488
rect 12069 3479 12127 3485
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13274 3519 13332 3525
rect 13274 3516 13286 3519
rect 13044 3488 13286 3516
rect 13044 3476 13050 3488
rect 13274 3485 13286 3488
rect 13320 3485 13332 3519
rect 13274 3479 13332 3485
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 16206 3516 16212 3528
rect 13955 3488 16212 3516
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3516 17463 3519
rect 18156 3516 18184 3556
rect 18782 3544 18788 3556
rect 18840 3544 18846 3596
rect 17451 3488 18184 3516
rect 18509 3519 18567 3525
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 18509 3485 18521 3519
rect 18555 3516 18567 3519
rect 18966 3516 18972 3528
rect 18555 3488 18972 3516
rect 18555 3485 18567 3488
rect 18509 3479 18567 3485
rect 11134 3420 11836 3448
rect 11900 3420 12296 3448
rect 11134 3417 11146 3420
rect 11088 3411 11146 3417
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8812 3352 8953 3380
rect 8812 3340 8818 3352
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 8941 3343 8999 3349
rect 9217 3383 9275 3389
rect 9217 3349 9229 3383
rect 9263 3349 9275 3383
rect 9766 3380 9772 3392
rect 9727 3352 9772 3380
rect 9217 3343 9275 3349
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 10870 3340 10876 3392
rect 10928 3380 10934 3392
rect 11790 3380 11796 3392
rect 10928 3352 11796 3380
rect 10928 3340 10934 3352
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 11900 3389 11928 3420
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3349 11943 3383
rect 12268 3380 12296 3420
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 13078 3448 13084 3460
rect 12400 3420 13084 3448
rect 12400 3408 12406 3420
rect 13078 3408 13084 3420
rect 13136 3408 13142 3460
rect 13446 3408 13452 3460
rect 13504 3448 13510 3460
rect 15228 3451 15286 3457
rect 13504 3420 14228 3448
rect 13504 3408 13510 3420
rect 12710 3380 12716 3392
rect 12268 3352 12716 3380
rect 11885 3343 11943 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 13725 3383 13783 3389
rect 13725 3380 13737 3383
rect 12860 3352 13737 3380
rect 12860 3340 12866 3352
rect 13725 3349 13737 3352
rect 13771 3349 13783 3383
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 13725 3343 13783 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 14200 3380 14228 3420
rect 15228 3417 15240 3451
rect 15274 3448 15286 3451
rect 15378 3448 15384 3460
rect 15274 3420 15384 3448
rect 15274 3417 15286 3420
rect 15228 3411 15286 3417
rect 15378 3408 15384 3420
rect 15436 3408 15442 3460
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 15810 3451 15868 3457
rect 15810 3448 15822 3451
rect 15620 3420 15822 3448
rect 15620 3408 15626 3420
rect 15810 3417 15822 3420
rect 15856 3417 15868 3451
rect 15810 3411 15868 3417
rect 17865 3451 17923 3457
rect 17865 3417 17877 3451
rect 17911 3448 17923 3451
rect 17954 3448 17960 3460
rect 17911 3420 17960 3448
rect 17911 3417 17923 3420
rect 17865 3411 17923 3417
rect 17954 3408 17960 3420
rect 18012 3448 18018 3460
rect 18524 3448 18552 3479
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 18012 3420 18552 3448
rect 18012 3408 18018 3420
rect 17770 3380 17776 3392
rect 14200 3352 17776 3380
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3881 3179 3939 3185
rect 3881 3145 3893 3179
rect 3927 3176 3939 3179
rect 4246 3176 4252 3188
rect 3927 3148 4108 3176
rect 4207 3148 4252 3176
rect 3927 3145 3939 3148
rect 3881 3139 3939 3145
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2774 3108 2780 3120
rect 1903 3080 2780 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 4080 3108 4108 3148
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 4801 3179 4859 3185
rect 4801 3176 4813 3179
rect 4672 3148 4813 3176
rect 4672 3136 4678 3148
rect 4801 3145 4813 3148
rect 4847 3145 4859 3179
rect 4801 3139 4859 3145
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 9306 3176 9312 3188
rect 5132 3148 9312 3176
rect 5132 3136 5138 3148
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 9824 3148 11560 3176
rect 9824 3136 9830 3148
rect 5810 3108 5816 3120
rect 2884 3080 3832 3108
rect 4080 3080 5816 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 1670 3040 1676 3052
rect 1627 3012 1676 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 2130 3040 2136 3052
rect 2091 3012 2136 3040
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2884 3049 2912 3080
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2869 3043 2927 3049
rect 2547 3012 2774 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2746 2972 2774 3012
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3326 3040 3332 3052
rect 3191 3012 3332 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 3694 3040 3700 3052
rect 3476 3012 3521 3040
rect 3655 3012 3700 3040
rect 3476 3000 3482 3012
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3804 3040 3832 3080
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 8202 3108 8208 3120
rect 6236 3080 8208 3108
rect 6236 3068 6242 3080
rect 4341 3043 4399 3049
rect 3804 3012 4108 3040
rect 3878 2972 3884 2984
rect 2746 2944 3884 2972
rect 3878 2932 3884 2944
rect 3936 2932 3942 2984
rect 2958 2864 2964 2916
rect 3016 2904 3022 2916
rect 3329 2907 3387 2913
rect 3329 2904 3341 2907
rect 3016 2876 3341 2904
rect 3016 2864 3022 2876
rect 3329 2873 3341 2876
rect 3375 2873 3387 2907
rect 3970 2904 3976 2916
rect 3329 2867 3387 2873
rect 3528 2876 3976 2904
rect 1394 2836 1400 2848
rect 1355 2808 1400 2836
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 1728 2808 2329 2836
rect 1728 2796 1734 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 2317 2799 2375 2805
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3528 2836 3556 2876
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4080 2904 4108 3012
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4387 3012 4752 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4614 2972 4620 2984
rect 4203 2944 4620 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 4724 2972 4752 3012
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5925 3043 5983 3049
rect 5925 3040 5937 3043
rect 4856 3012 5937 3040
rect 4856 3000 4862 3012
rect 5925 3009 5937 3012
rect 5971 3040 5983 3043
rect 6086 3040 6092 3052
rect 5971 3012 6092 3040
rect 5971 3009 5983 3012
rect 5925 3003 5983 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7852 3049 7880 3080
rect 8202 3068 8208 3080
rect 8260 3108 8266 3120
rect 11330 3108 11336 3120
rect 8260 3080 11336 3108
rect 8260 3068 8266 3080
rect 7581 3043 7639 3049
rect 7581 3040 7593 3043
rect 7156 3012 7593 3040
rect 7156 3000 7162 3012
rect 7581 3009 7593 3012
rect 7627 3040 7639 3043
rect 7837 3043 7895 3049
rect 7627 3012 7788 3040
rect 7627 3009 7639 3012
rect 7581 3003 7639 3009
rect 5166 2972 5172 2984
rect 4724 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6178 2972 6184 2984
rect 6139 2944 6184 2972
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 7760 2972 7788 3012
rect 7837 3009 7849 3043
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 8021 2975 8079 2981
rect 7760 2944 7880 2972
rect 4982 2904 4988 2916
rect 4080 2876 4988 2904
rect 4982 2864 4988 2876
rect 5040 2864 5046 2916
rect 7852 2904 7880 2944
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8110 2972 8116 2984
rect 8067 2944 8116 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8220 2972 8248 3068
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8444 3012 8489 3040
rect 8444 3000 8450 3012
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 9968 3049 9996 3080
rect 11330 3068 11336 3080
rect 11388 3068 11394 3120
rect 8737 3043 8795 3049
rect 8737 3040 8749 3043
rect 8628 3012 8749 3040
rect 8628 3000 8634 3012
rect 8737 3009 8749 3012
rect 8783 3009 8795 3043
rect 8737 3003 8795 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 10226 3049 10232 3052
rect 10220 3040 10232 3049
rect 10100 3012 10232 3040
rect 10100 3000 10106 3012
rect 10220 3003 10232 3012
rect 10226 3000 10232 3003
rect 10284 3000 10290 3052
rect 11532 3049 11560 3148
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 11977 3179 12035 3185
rect 11977 3176 11989 3179
rect 11848 3148 11989 3176
rect 11848 3136 11854 3148
rect 11977 3145 11989 3148
rect 12023 3145 12035 3179
rect 11977 3139 12035 3145
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13446 3176 13452 3188
rect 12492 3148 13452 3176
rect 12492 3136 12498 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 14844 3148 15608 3176
rect 13112 3111 13170 3117
rect 13112 3077 13124 3111
rect 13158 3108 13170 3111
rect 13722 3108 13728 3120
rect 13158 3080 13728 3108
rect 13158 3077 13170 3080
rect 13112 3071 13170 3077
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 13814 3068 13820 3120
rect 13872 3108 13878 3120
rect 14584 3111 14642 3117
rect 14584 3108 14596 3111
rect 13872 3080 14596 3108
rect 13872 3068 13878 3080
rect 14584 3077 14596 3080
rect 14630 3108 14642 3111
rect 14844 3108 14872 3148
rect 15470 3108 15476 3120
rect 14630 3080 14872 3108
rect 14936 3080 15476 3108
rect 14630 3077 14642 3080
rect 14584 3071 14642 3077
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13320 3012 13369 3040
rect 13320 3000 13326 3012
rect 13357 3009 13369 3012
rect 13403 3040 13415 3043
rect 13538 3040 13544 3052
rect 13403 3012 13544 3040
rect 13403 3009 13415 3012
rect 13357 3003 13415 3009
rect 13538 3000 13544 3012
rect 13596 3040 13602 3052
rect 14936 3049 14964 3080
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15580 3108 15608 3148
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 16080 3148 16313 3176
rect 16080 3136 16086 3148
rect 16301 3145 16313 3148
rect 16347 3145 16359 3179
rect 16301 3139 16359 3145
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 16908 3148 16957 3176
rect 16908 3136 16914 3148
rect 16945 3145 16957 3148
rect 16991 3145 17003 3179
rect 16945 3139 17003 3145
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17184 3148 17325 3176
rect 17184 3136 17190 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17451 3148 17785 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 18506 3176 18512 3188
rect 18187 3148 18512 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 15580 3080 18368 3108
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 13596 3012 14841 3040
rect 13596 3000 13602 3012
rect 14829 3009 14841 3012
rect 14875 3040 14887 3043
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14875 3012 14933 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15188 3043 15246 3049
rect 15188 3009 15200 3043
rect 15234 3040 15246 3043
rect 15562 3040 15568 3052
rect 15234 3012 15568 3040
rect 15234 3009 15246 3012
rect 15188 3003 15246 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16448 3012 16865 3040
rect 16448 3000 16454 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 17644 3012 18245 3040
rect 17644 3000 17650 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 8294 2972 8300 2984
rect 8220 2944 8300 2972
rect 8294 2932 8300 2944
rect 8352 2972 8358 2984
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8352 2944 8493 2972
rect 8352 2932 8358 2944
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 17497 2975 17555 2981
rect 8481 2935 8539 2941
rect 10980 2944 11836 2972
rect 7852 2876 8156 2904
rect 8128 2848 8156 2876
rect 2832 2808 3556 2836
rect 2832 2796 2838 2808
rect 3602 2796 3608 2848
rect 3660 2836 3666 2848
rect 4706 2836 4712 2848
rect 3660 2808 3705 2836
rect 4667 2808 4712 2836
rect 3660 2796 3666 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 6457 2839 6515 2845
rect 6457 2805 6469 2839
rect 6503 2836 6515 2839
rect 7190 2836 7196 2848
rect 6503 2808 7196 2836
rect 6503 2805 6515 2808
rect 6457 2799 6515 2805
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 8110 2796 8116 2848
rect 8168 2796 8174 2848
rect 8205 2839 8263 2845
rect 8205 2805 8217 2839
rect 8251 2836 8263 2839
rect 8662 2836 8668 2848
rect 8251 2808 8668 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 9674 2836 9680 2848
rect 9272 2808 9680 2836
rect 9272 2796 9278 2808
rect 9674 2796 9680 2808
rect 9732 2836 9738 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9732 2808 9873 2836
rect 9732 2796 9738 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10980 2836 11008 2944
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 11204 2876 11713 2904
rect 11204 2864 11210 2876
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 11808 2904 11836 2944
rect 17497 2941 17509 2975
rect 17543 2972 17555 2975
rect 17770 2972 17776 2984
rect 17543 2944 17776 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18340 2981 18368 3080
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 16485 2907 16543 2913
rect 11808 2876 12434 2904
rect 11701 2867 11759 2873
rect 10376 2808 11008 2836
rect 11333 2839 11391 2845
rect 10376 2796 10382 2808
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 11422 2836 11428 2848
rect 11379 2808 11428 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 12406 2836 12434 2876
rect 16485 2873 16497 2907
rect 16531 2904 16543 2907
rect 17954 2904 17960 2916
rect 16531 2876 17960 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 17954 2864 17960 2876
rect 18012 2864 18018 2916
rect 13170 2836 13176 2848
rect 12406 2808 13176 2836
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13630 2796 13636 2848
rect 13688 2836 13694 2848
rect 15562 2836 15568 2848
rect 13688 2808 15568 2836
rect 13688 2796 13694 2808
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 16850 2836 16856 2848
rect 16715 2808 16856 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 3878 2632 3884 2644
rect 3839 2604 3884 2632
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 5258 2632 5264 2644
rect 4203 2604 5264 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 9122 2632 9128 2644
rect 5951 2604 8432 2632
rect 9083 2604 9128 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 1210 2524 1216 2576
rect 1268 2564 1274 2576
rect 2593 2567 2651 2573
rect 2593 2564 2605 2567
rect 1268 2536 2605 2564
rect 1268 2524 1274 2536
rect 2593 2533 2605 2536
rect 2639 2533 2651 2567
rect 3694 2564 3700 2576
rect 2593 2527 2651 2533
rect 3160 2536 3700 2564
rect 2866 2496 2872 2508
rect 2424 2468 2872 2496
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2314 2428 2320 2440
rect 2087 2400 2320 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2424 2437 2452 2468
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3160 2428 3188 2536
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 6181 2567 6239 2573
rect 4764 2536 5488 2564
rect 4764 2524 4770 2536
rect 4062 2496 4068 2508
rect 3252 2468 4068 2496
rect 3252 2437 3280 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2496 4675 2499
rect 4982 2496 4988 2508
rect 4663 2468 4988 2496
rect 4663 2465 4675 2468
rect 4617 2459 4675 2465
rect 2823 2400 3188 2428
rect 3237 2431 3295 2437
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3344 2360 3372 2391
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3660 2400 3985 2428
rect 3660 2388 3666 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 3016 2332 3372 2360
rect 4540 2360 4568 2459
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 5460 2505 5488 2536
rect 6181 2533 6193 2567
rect 6227 2533 6239 2567
rect 6181 2527 6239 2533
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 5445 2499 5503 2505
rect 5445 2465 5457 2499
rect 5491 2465 5503 2499
rect 6196 2496 6224 2527
rect 8404 2496 8432 2604
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 11514 2632 11520 2644
rect 9640 2604 9812 2632
rect 11475 2604 11520 2632
rect 9640 2592 9646 2604
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 9490 2564 9496 2576
rect 8619 2536 9496 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 9784 2505 9812 2604
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11974 2592 11980 2644
rect 12032 2632 12038 2644
rect 13541 2635 13599 2641
rect 13541 2632 13553 2635
rect 12032 2604 13553 2632
rect 12032 2592 12038 2604
rect 13541 2601 13553 2604
rect 13587 2601 13599 2635
rect 13541 2595 13599 2601
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 16025 2635 16083 2641
rect 16025 2632 16037 2635
rect 14792 2604 16037 2632
rect 14792 2592 14798 2604
rect 16025 2601 16037 2604
rect 16071 2601 16083 2635
rect 16025 2595 16083 2601
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 16264 2604 16313 2632
rect 16264 2592 16270 2604
rect 16301 2601 16313 2604
rect 16347 2601 16359 2635
rect 16301 2595 16359 2601
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 17770 2632 17776 2644
rect 17267 2604 17776 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18414 2632 18420 2644
rect 18375 2604 18420 2632
rect 18414 2592 18420 2604
rect 18472 2592 18478 2644
rect 13170 2564 13176 2576
rect 13131 2536 13176 2564
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 15562 2524 15568 2576
rect 15620 2564 15626 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 15620 2536 15761 2564
rect 15620 2524 15626 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 15749 2527 15807 2533
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 6196 2468 6684 2496
rect 8404 2468 9597 2496
rect 5445 2459 5503 2465
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 4798 2428 4804 2440
rect 4755 2400 4804 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 5368 2428 5396 2459
rect 5994 2428 6000 2440
rect 5368 2400 5856 2428
rect 5955 2400 6000 2428
rect 4614 2360 4620 2372
rect 4540 2332 4620 2360
rect 3016 2320 3022 2332
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 5537 2363 5595 2369
rect 5537 2360 5549 2363
rect 5092 2332 5549 2360
rect 1854 2292 1860 2304
rect 1815 2264 1860 2292
rect 1854 2252 1860 2264
rect 1912 2252 1918 2304
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2096 2264 2237 2292
rect 2096 2252 2102 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 3053 2295 3111 2301
rect 3053 2292 3065 2295
rect 2924 2264 3065 2292
rect 2924 2252 2930 2264
rect 3053 2261 3065 2264
rect 3099 2261 3111 2295
rect 3053 2255 3111 2261
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3694 2292 3700 2304
rect 3559 2264 3700 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3694 2252 3700 2264
rect 3752 2252 3758 2304
rect 5092 2301 5120 2332
rect 5537 2329 5549 2332
rect 5583 2329 5595 2363
rect 5828 2360 5856 2400
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 6454 2428 6460 2440
rect 6411 2400 6460 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 6656 2437 6684 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 11330 2496 11336 2508
rect 9815 2468 10364 2496
rect 11291 2468 11336 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8352 2400 8401 2428
rect 8352 2388 8358 2400
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 8754 2428 8760 2440
rect 8715 2400 8760 2428
rect 8389 2391 8447 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2428 9091 2431
rect 10042 2428 10048 2440
rect 9079 2400 10048 2428
rect 9079 2397 9091 2400
rect 9033 2391 9091 2397
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10336 2428 10364 2468
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 13262 2496 13268 2508
rect 12943 2468 13268 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 14090 2496 14096 2508
rect 13464 2468 14096 2496
rect 12986 2428 12992 2440
rect 10336 2400 12434 2428
rect 12947 2400 12992 2428
rect 7282 2360 7288 2372
rect 5828 2332 7288 2360
rect 5537 2323 5595 2329
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2261 5135 2295
rect 6546 2292 6552 2304
rect 6507 2264 6552 2292
rect 5077 2255 5135 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 6825 2295 6883 2301
rect 6825 2261 6837 2295
rect 6871 2292 6883 2295
rect 6914 2292 6920 2304
rect 6871 2264 6920 2292
rect 6871 2261 6883 2264
rect 6825 2255 6883 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7024 2301 7052 2332
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7374 2320 7380 2372
rect 7432 2360 7438 2372
rect 8144 2363 8202 2369
rect 8144 2360 8156 2363
rect 7432 2332 8156 2360
rect 7432 2320 7438 2332
rect 8144 2329 8156 2332
rect 8190 2360 8202 2363
rect 9214 2360 9220 2372
rect 8190 2332 9220 2360
rect 8190 2329 8202 2332
rect 8144 2323 8202 2329
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 9398 2320 9404 2372
rect 9456 2360 9462 2372
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 9456 2332 9505 2360
rect 9456 2320 9462 2332
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 11066 2363 11124 2369
rect 11066 2360 11078 2363
rect 9493 2323 9551 2329
rect 9600 2332 11078 2360
rect 7009 2295 7067 2301
rect 7009 2261 7021 2295
rect 7055 2261 7067 2295
rect 7009 2255 7067 2261
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 9600 2292 9628 2332
rect 11066 2329 11078 2332
rect 11112 2360 11124 2363
rect 12406 2360 12434 2400
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 13136 2400 13369 2428
rect 13136 2388 13142 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 12630 2363 12688 2369
rect 12630 2360 12642 2363
rect 11112 2332 11192 2360
rect 12406 2332 12642 2360
rect 11112 2329 11124 2332
rect 11066 2323 11124 2329
rect 7984 2264 9628 2292
rect 7984 2252 7990 2264
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9824 2264 9965 2292
rect 9824 2252 9830 2264
rect 9953 2261 9965 2264
rect 9999 2292 10011 2295
rect 10686 2292 10692 2304
rect 9999 2264 10692 2292
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 11164 2292 11192 2332
rect 12630 2329 12642 2332
rect 12676 2329 12688 2363
rect 12630 2323 12688 2329
rect 13464 2292 13492 2468
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16850 2496 16856 2508
rect 16224 2468 16856 2496
rect 13722 2428 13728 2440
rect 13683 2400 13728 2428
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 16224 2437 16252 2468
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 13924 2400 15577 2428
rect 13924 2301 13952 2400
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 16209 2431 16267 2437
rect 16209 2397 16221 2431
rect 16255 2397 16267 2431
rect 16209 2391 16267 2397
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16356 2400 16497 2428
rect 16356 2388 16362 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 16761 2431 16819 2437
rect 16761 2397 16773 2431
rect 16807 2397 16819 2431
rect 17402 2428 17408 2440
rect 17363 2400 17408 2428
rect 16761 2391 16819 2397
rect 14642 2320 14648 2372
rect 14700 2360 14706 2372
rect 15206 2363 15264 2369
rect 15206 2360 15218 2363
rect 14700 2332 15218 2360
rect 14700 2320 14706 2332
rect 15206 2329 15218 2332
rect 15252 2329 15264 2363
rect 15206 2323 15264 2329
rect 11164 2264 13492 2292
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2261 13967 2295
rect 14090 2292 14096 2304
rect 14051 2264 14096 2292
rect 13909 2255 13967 2261
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 16776 2292 16804 2391
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 17494 2388 17500 2440
rect 17552 2428 17558 2440
rect 17862 2428 17868 2440
rect 17552 2400 17597 2428
rect 17823 2400 17868 2428
rect 17552 2388 17558 2400
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18233 2431 18291 2437
rect 18233 2428 18245 2431
rect 18196 2400 18245 2428
rect 18196 2388 18202 2400
rect 18233 2397 18245 2400
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 16942 2292 16948 2304
rect 14884 2264 16804 2292
rect 16903 2264 16948 2292
rect 14884 2252 14890 2264
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17770 2292 17776 2304
rect 17727 2264 17776 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 1486 2048 1492 2100
rect 1544 2088 1550 2100
rect 1544 2060 2774 2088
rect 1544 2048 1550 2060
rect 2746 1884 2774 2060
rect 4614 2048 4620 2100
rect 4672 2088 4678 2100
rect 7374 2088 7380 2100
rect 4672 2060 7380 2088
rect 4672 2048 4678 2060
rect 7374 2048 7380 2060
rect 7432 2048 7438 2100
rect 14182 2048 14188 2100
rect 14240 2088 14246 2100
rect 17862 2088 17868 2100
rect 14240 2060 17868 2088
rect 14240 2048 14246 2060
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 6546 1980 6552 2032
rect 6604 2020 6610 2032
rect 12986 2020 12992 2032
rect 6604 1992 12992 2020
rect 6604 1980 6610 1992
rect 12986 1980 12992 1992
rect 13044 1980 13050 2032
rect 13354 1980 13360 2032
rect 13412 2020 13418 2032
rect 16942 2020 16948 2032
rect 13412 1992 16948 2020
rect 13412 1980 13418 1992
rect 16942 1980 16948 1992
rect 17000 1980 17006 2032
rect 3050 1912 3056 1964
rect 3108 1952 3114 1964
rect 7926 1952 7932 1964
rect 3108 1924 7932 1952
rect 3108 1912 3114 1924
rect 7926 1912 7932 1924
rect 7984 1912 7990 1964
rect 8110 1912 8116 1964
rect 8168 1952 8174 1964
rect 14090 1952 14096 1964
rect 8168 1924 14096 1952
rect 8168 1912 8174 1924
rect 14090 1912 14096 1924
rect 14148 1912 14154 1964
rect 9766 1884 9772 1896
rect 2746 1856 9772 1884
rect 9766 1844 9772 1856
rect 9824 1844 9830 1896
rect 12710 1776 12716 1828
rect 12768 1816 12774 1828
rect 15378 1816 15384 1828
rect 12768 1788 15384 1816
rect 12768 1776 12774 1788
rect 15378 1776 15384 1788
rect 15436 1776 15442 1828
<< via1 >>
rect 2320 14968 2372 15020
rect 6552 14968 6604 15020
rect 5908 14900 5960 14952
rect 15292 14900 15344 14952
rect 3608 14832 3660 14884
rect 6920 14832 6972 14884
rect 4436 14764 4488 14816
rect 5448 14764 5500 14816
rect 15200 14764 15252 14816
rect 16212 14764 16264 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 2780 14560 2832 14612
rect 5724 14603 5776 14612
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 2780 14424 2832 14476
rect 3516 14424 3568 14476
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2964 14356 3016 14408
rect 4068 14356 4120 14408
rect 4252 14356 4304 14408
rect 4436 14356 4488 14408
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 6552 14603 6604 14612
rect 6552 14569 6561 14603
rect 6561 14569 6595 14603
rect 6595 14569 6604 14603
rect 6552 14560 6604 14569
rect 7472 14560 7524 14612
rect 10140 14603 10192 14612
rect 5540 14492 5592 14544
rect 3056 14288 3108 14340
rect 5540 14356 5592 14408
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 11980 14560 12032 14612
rect 14556 14603 14608 14612
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 15476 14492 15528 14544
rect 15200 14424 15252 14476
rect 15660 14424 15712 14476
rect 10876 14356 10928 14408
rect 12808 14356 12860 14408
rect 13820 14356 13872 14408
rect 15384 14356 15436 14408
rect 16856 14424 16908 14476
rect 16396 14399 16448 14408
rect 8116 14288 8168 14340
rect 15200 14288 15252 14340
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 16028 14331 16080 14340
rect 16028 14297 16037 14331
rect 16037 14297 16071 14331
rect 16071 14297 16080 14331
rect 16028 14288 16080 14297
rect 16212 14288 16264 14340
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 17868 14356 17920 14408
rect 3148 14220 3200 14272
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 4896 14263 4948 14272
rect 4896 14229 4905 14263
rect 4905 14229 4939 14263
rect 4939 14229 4948 14263
rect 4896 14220 4948 14229
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 5264 14220 5316 14272
rect 5448 14220 5500 14272
rect 10232 14220 10284 14272
rect 14096 14220 14148 14272
rect 16120 14220 16172 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 4436 14016 4488 14068
rect 5264 14016 5316 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6920 14059 6972 14068
rect 6920 14025 6929 14059
rect 6929 14025 6963 14059
rect 6963 14025 6972 14059
rect 6920 14016 6972 14025
rect 12808 14059 12860 14068
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 2780 13880 2832 13932
rect 2964 13880 3016 13932
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 4068 13880 4120 13932
rect 1768 13812 1820 13864
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 3424 13812 3476 13864
rect 3608 13812 3660 13864
rect 3792 13812 3844 13864
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 4712 13855 4764 13864
rect 4712 13821 4721 13855
rect 4721 13821 4755 13855
rect 4755 13821 4764 13855
rect 4712 13812 4764 13821
rect 4988 13812 5040 13864
rect 5080 13812 5132 13864
rect 6000 13812 6052 13864
rect 8944 13812 8996 13864
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 12900 13880 12952 13932
rect 13820 13880 13872 13932
rect 15660 13948 15712 14000
rect 17132 13991 17184 14000
rect 17132 13957 17141 13991
rect 17141 13957 17175 13991
rect 17175 13957 17184 13991
rect 17132 13948 17184 13957
rect 17500 13991 17552 14000
rect 17500 13957 17509 13991
rect 17509 13957 17543 13991
rect 17543 13957 17552 13991
rect 17500 13948 17552 13957
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16028 13880 16080 13932
rect 16304 13880 16356 13932
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 13544 13855 13596 13864
rect 13544 13821 13553 13855
rect 13553 13821 13587 13855
rect 13587 13821 13596 13855
rect 13544 13812 13596 13821
rect 14004 13812 14056 13864
rect 1124 13744 1176 13796
rect 3056 13676 3108 13728
rect 4068 13744 4120 13796
rect 3884 13676 3936 13728
rect 4896 13676 4948 13728
rect 15292 13787 15344 13796
rect 15292 13753 15301 13787
rect 15301 13753 15335 13787
rect 15335 13753 15344 13787
rect 15292 13744 15344 13753
rect 16120 13744 16172 13796
rect 6460 13676 6512 13728
rect 10876 13676 10928 13728
rect 15200 13676 15252 13728
rect 15660 13676 15712 13728
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 18328 13812 18380 13864
rect 16856 13787 16908 13796
rect 16856 13753 16865 13787
rect 16865 13753 16899 13787
rect 16899 13753 16908 13787
rect 16856 13744 16908 13753
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 3056 13472 3108 13524
rect 3424 13472 3476 13524
rect 4620 13472 4672 13524
rect 6276 13472 6328 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 16764 13404 16816 13456
rect 17776 13404 17828 13456
rect 3056 13379 3108 13388
rect 3056 13345 3065 13379
rect 3065 13345 3099 13379
rect 3099 13345 3108 13379
rect 3056 13336 3108 13345
rect 3884 13336 3936 13388
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 3424 13268 3476 13320
rect 4712 13268 4764 13320
rect 6092 13336 6144 13388
rect 6920 13336 6972 13388
rect 17960 13379 18012 13388
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 6552 13268 6604 13320
rect 6828 13268 6880 13320
rect 15108 13311 15160 13320
rect 2872 13200 2924 13252
rect 3700 13200 3752 13252
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 5816 13243 5868 13252
rect 5816 13209 5825 13243
rect 5825 13209 5859 13243
rect 5859 13209 5868 13243
rect 5816 13200 5868 13209
rect 6000 13200 6052 13252
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 13268 13200 13320 13252
rect 15384 13200 15436 13252
rect 1216 13132 1268 13184
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 2964 13132 3016 13184
rect 3976 13175 4028 13184
rect 3976 13141 3985 13175
rect 3985 13141 4019 13175
rect 4019 13141 4028 13175
rect 3976 13132 4028 13141
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4988 13175 5040 13184
rect 4528 13132 4580 13141
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5080 13132 5132 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 11152 13132 11204 13184
rect 14832 13132 14884 13184
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 17500 13243 17552 13252
rect 17224 13175 17276 13184
rect 17224 13141 17233 13175
rect 17233 13141 17267 13175
rect 17267 13141 17276 13175
rect 17224 13132 17276 13141
rect 17500 13209 17509 13243
rect 17509 13209 17543 13243
rect 17543 13209 17552 13243
rect 17500 13200 17552 13209
rect 18788 13132 18840 13184
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2136 12928 2188 12980
rect 3056 12928 3108 12980
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 5080 12928 5132 12980
rect 6828 12928 6880 12980
rect 7380 12928 7432 12980
rect 17592 12928 17644 12980
rect 6460 12860 6512 12912
rect 7012 12860 7064 12912
rect 2504 12792 2556 12844
rect 4896 12792 4948 12844
rect 5632 12792 5684 12844
rect 13452 12903 13504 12912
rect 13452 12869 13461 12903
rect 13461 12869 13495 12903
rect 13495 12869 13504 12903
rect 13452 12860 13504 12869
rect 17500 12860 17552 12912
rect 10600 12792 10652 12844
rect 12624 12792 12676 12844
rect 16304 12835 16356 12844
rect 16304 12801 16313 12835
rect 16313 12801 16347 12835
rect 16347 12801 16356 12835
rect 16304 12792 16356 12801
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 17316 12792 17368 12844
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 4528 12724 4580 12776
rect 2780 12656 2832 12708
rect 2964 12656 3016 12708
rect 3976 12656 4028 12708
rect 6368 12724 6420 12776
rect 7380 12724 7432 12776
rect 7472 12724 7524 12776
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 14648 12724 14700 12776
rect 17684 12767 17736 12776
rect 17684 12733 17693 12767
rect 17693 12733 17727 12767
rect 17727 12733 17736 12767
rect 17684 12724 17736 12733
rect 6092 12656 6144 12708
rect 9220 12656 9272 12708
rect 16120 12656 16172 12708
rect 3516 12588 3568 12640
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 6000 12588 6052 12640
rect 6736 12588 6788 12640
rect 6828 12588 6880 12640
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 13728 12588 13780 12640
rect 16396 12631 16448 12640
rect 16396 12597 16405 12631
rect 16405 12597 16439 12631
rect 16439 12597 16448 12631
rect 16396 12588 16448 12597
rect 17040 12588 17092 12640
rect 17500 12588 17552 12640
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 18144 12588 18196 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2872 12384 2924 12436
rect 4252 12384 4304 12436
rect 5080 12384 5132 12436
rect 9680 12384 9732 12436
rect 10232 12316 10284 12368
rect 12532 12384 12584 12436
rect 13452 12384 13504 12436
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 10416 12316 10468 12368
rect 12440 12316 12492 12368
rect 14096 12316 14148 12368
rect 14832 12316 14884 12368
rect 3516 12291 3568 12300
rect 3516 12257 3525 12291
rect 3525 12257 3559 12291
rect 3559 12257 3568 12291
rect 3516 12248 3568 12257
rect 3700 12248 3752 12300
rect 4528 12248 4580 12300
rect 4896 12291 4948 12300
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 2044 12112 2096 12164
rect 2688 12180 2740 12232
rect 4160 12180 4212 12232
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 5080 12180 5132 12232
rect 5632 12180 5684 12232
rect 7380 12248 7432 12300
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 7288 12180 7340 12232
rect 10968 12248 11020 12300
rect 12072 12248 12124 12300
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 17868 12384 17920 12436
rect 17960 12316 18012 12368
rect 14648 12248 14700 12257
rect 8116 12180 8168 12232
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 9772 12180 9824 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 12992 12180 13044 12232
rect 13912 12180 13964 12232
rect 14004 12180 14056 12232
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 17592 12248 17644 12300
rect 14556 12180 14608 12189
rect 2780 12087 2832 12096
rect 2780 12053 2789 12087
rect 2789 12053 2823 12087
rect 2823 12053 2832 12087
rect 2780 12044 2832 12053
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 4068 12044 4120 12096
rect 4804 12044 4856 12096
rect 5264 12044 5316 12096
rect 5724 12044 5776 12096
rect 5816 12044 5868 12096
rect 7012 12044 7064 12096
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 10416 12112 10468 12164
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 8484 12044 8536 12096
rect 9220 12044 9272 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12624 12044 12676 12096
rect 13360 12044 13412 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 14004 12044 14056 12096
rect 14188 12112 14240 12164
rect 17684 12223 17736 12232
rect 16120 12112 16172 12164
rect 16488 12155 16540 12164
rect 16488 12121 16497 12155
rect 16497 12121 16531 12155
rect 16531 12121 16540 12155
rect 16488 12112 16540 12121
rect 15936 12087 15988 12096
rect 15936 12053 15945 12087
rect 15945 12053 15979 12087
rect 15979 12053 15988 12087
rect 15936 12044 15988 12053
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 16304 12044 16356 12096
rect 17132 12044 17184 12096
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 17776 12044 17828 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 3884 11840 3936 11892
rect 4068 11883 4120 11892
rect 4068 11849 4077 11883
rect 4077 11849 4111 11883
rect 4111 11849 4120 11883
rect 4068 11840 4120 11849
rect 5080 11840 5132 11892
rect 5264 11840 5316 11892
rect 5724 11840 5776 11892
rect 6276 11840 6328 11892
rect 7104 11840 7156 11892
rect 7656 11840 7708 11892
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 8484 11883 8536 11892
rect 7748 11840 7800 11849
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 9772 11840 9824 11892
rect 11980 11840 12032 11892
rect 4988 11772 5040 11824
rect 5816 11772 5868 11824
rect 9220 11772 9272 11824
rect 9496 11772 9548 11824
rect 9680 11772 9732 11824
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 1676 11704 1728 11756
rect 1124 11500 1176 11552
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 2136 11568 2188 11620
rect 2504 11611 2556 11620
rect 2504 11577 2513 11611
rect 2513 11577 2547 11611
rect 2547 11577 2556 11611
rect 2504 11568 2556 11577
rect 2780 11636 2832 11688
rect 4160 11704 4212 11756
rect 3516 11636 3568 11688
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 7104 11704 7156 11756
rect 9312 11747 9364 11756
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 6092 11636 6144 11688
rect 6736 11636 6788 11688
rect 4160 11568 4212 11620
rect 4252 11568 4304 11620
rect 6552 11568 6604 11620
rect 6920 11568 6972 11620
rect 7104 11568 7156 11620
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 7748 11568 7800 11620
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9588 11704 9640 11756
rect 12440 11772 12492 11824
rect 14188 11772 14240 11824
rect 14556 11772 14608 11824
rect 13452 11747 13504 11756
rect 9220 11636 9272 11688
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 10140 11636 10192 11688
rect 3516 11500 3568 11552
rect 4068 11500 4120 11552
rect 5080 11500 5132 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6368 11500 6420 11552
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7932 11500 7984 11552
rect 8392 11500 8444 11552
rect 9312 11500 9364 11552
rect 10416 11568 10468 11620
rect 10968 11679 11020 11688
rect 10968 11645 10977 11679
rect 10977 11645 11011 11679
rect 11011 11645 11020 11679
rect 10968 11636 11020 11645
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 11980 11636 12032 11645
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12716 11636 12768 11688
rect 13636 11704 13688 11756
rect 14924 11704 14976 11756
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 16856 11704 16908 11756
rect 17224 11772 17276 11824
rect 17500 11704 17552 11756
rect 18052 11747 18104 11756
rect 18052 11713 18061 11747
rect 18061 11713 18095 11747
rect 18095 11713 18104 11747
rect 18052 11704 18104 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 11244 11568 11296 11620
rect 14556 11611 14608 11620
rect 14556 11577 14565 11611
rect 14565 11577 14599 11611
rect 14599 11577 14608 11611
rect 14556 11568 14608 11577
rect 16212 11636 16264 11688
rect 16488 11636 16540 11688
rect 17132 11636 17184 11688
rect 15844 11568 15896 11620
rect 9864 11500 9916 11552
rect 10508 11500 10560 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 14372 11500 14424 11552
rect 14740 11543 14792 11552
rect 14740 11509 14749 11543
rect 14749 11509 14783 11543
rect 14783 11509 14792 11543
rect 14740 11500 14792 11509
rect 15476 11500 15528 11552
rect 15752 11500 15804 11552
rect 18696 11568 18748 11620
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 16120 11500 16172 11509
rect 16396 11500 16448 11552
rect 16948 11500 17000 11552
rect 17868 11500 17920 11552
rect 18236 11500 18288 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 1768 11296 1820 11348
rect 3792 11296 3844 11348
rect 1860 11228 1912 11280
rect 2412 11160 2464 11212
rect 4160 11228 4212 11280
rect 4804 11296 4856 11348
rect 6644 11296 6696 11348
rect 7564 11296 7616 11348
rect 8576 11296 8628 11348
rect 11060 11296 11112 11348
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 15384 11296 15436 11348
rect 16396 11296 16448 11348
rect 16856 11339 16908 11348
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 4252 11160 4304 11212
rect 4896 11228 4948 11280
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6276 11160 6328 11212
rect 7472 11228 7524 11280
rect 2688 11024 2740 11076
rect 3976 11024 4028 11076
rect 7012 11160 7064 11212
rect 7656 11160 7708 11212
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 7564 11135 7616 11144
rect 6828 11092 6880 11101
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 6552 11024 6604 11076
rect 6920 11024 6972 11076
rect 7288 11024 7340 11076
rect 8576 11160 8628 11212
rect 10416 11228 10468 11280
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 3148 10956 3200 11008
rect 4252 10956 4304 11008
rect 4988 10956 5040 11008
rect 5264 10956 5316 11008
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 8484 11024 8536 11076
rect 9588 11092 9640 11144
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 8760 11024 8812 11076
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 10600 10956 10652 11008
rect 11244 11160 11296 11212
rect 14924 11228 14976 11280
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 18972 11228 19024 11280
rect 11520 11024 11572 11076
rect 13452 11160 13504 11212
rect 13728 11160 13780 11212
rect 15568 11160 15620 11212
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 15936 11160 15988 11212
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13176 11092 13228 11144
rect 14372 11092 14424 11144
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 16212 11135 16264 11144
rect 16212 11101 16221 11135
rect 16221 11101 16255 11135
rect 16255 11101 16264 11135
rect 16212 11092 16264 11101
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 16580 11092 16632 11144
rect 17132 11160 17184 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 17684 11135 17736 11144
rect 13728 11024 13780 11076
rect 13820 11067 13872 11076
rect 13820 11033 13829 11067
rect 13829 11033 13863 11067
rect 13863 11033 13872 11067
rect 13820 11024 13872 11033
rect 16672 11024 16724 11076
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 17408 11024 17460 11076
rect 10968 10956 11020 11008
rect 11796 10956 11848 11008
rect 13452 10999 13504 11008
rect 13452 10965 13461 10999
rect 13461 10965 13495 10999
rect 13495 10965 13504 10999
rect 13452 10956 13504 10965
rect 15108 10999 15160 11008
rect 15108 10965 15117 10999
rect 15117 10965 15151 10999
rect 15151 10965 15160 10999
rect 15108 10956 15160 10965
rect 15936 10956 15988 11008
rect 17040 10956 17092 11008
rect 17224 10999 17276 11008
rect 17224 10965 17233 10999
rect 17233 10965 17267 10999
rect 17267 10965 17276 10999
rect 17224 10956 17276 10965
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 1952 10752 2004 10804
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 2228 10684 2280 10736
rect 3976 10752 4028 10804
rect 4528 10752 4580 10804
rect 4988 10752 5040 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 6368 10752 6420 10804
rect 2320 10616 2372 10668
rect 2688 10616 2740 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 3516 10548 3568 10600
rect 4988 10616 5040 10668
rect 5172 10616 5224 10668
rect 5816 10616 5868 10668
rect 6184 10616 6236 10668
rect 8852 10752 8904 10804
rect 10232 10752 10284 10804
rect 12624 10752 12676 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 13452 10752 13504 10804
rect 15108 10752 15160 10804
rect 15200 10795 15252 10804
rect 15200 10761 15209 10795
rect 15209 10761 15243 10795
rect 15243 10761 15252 10795
rect 15200 10752 15252 10761
rect 11980 10684 12032 10736
rect 3056 10480 3108 10532
rect 4528 10480 4580 10532
rect 5080 10548 5132 10600
rect 5632 10548 5684 10600
rect 6460 10548 6512 10600
rect 9772 10616 9824 10668
rect 10968 10616 11020 10668
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 13636 10684 13688 10736
rect 13820 10684 13872 10736
rect 14740 10684 14792 10736
rect 14188 10616 14240 10668
rect 16120 10752 16172 10804
rect 16672 10795 16724 10804
rect 16672 10761 16681 10795
rect 16681 10761 16715 10795
rect 16715 10761 16724 10795
rect 16672 10752 16724 10761
rect 15844 10684 15896 10736
rect 6828 10548 6880 10600
rect 7012 10548 7064 10600
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 4344 10412 4396 10464
rect 8024 10480 8076 10532
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 6000 10412 6052 10464
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7472 10412 7524 10464
rect 8208 10412 8260 10464
rect 8576 10548 8628 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 10416 10548 10468 10600
rect 11612 10548 11664 10600
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 13452 10591 13504 10600
rect 12440 10548 12492 10557
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 13820 10548 13872 10600
rect 14648 10548 14700 10600
rect 15476 10548 15528 10600
rect 8944 10412 8996 10464
rect 10232 10412 10284 10464
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 12808 10480 12860 10532
rect 13176 10480 13228 10532
rect 16764 10616 16816 10668
rect 17224 10752 17276 10804
rect 11796 10412 11848 10464
rect 11980 10412 12032 10464
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 14464 10412 14516 10464
rect 15200 10412 15252 10464
rect 16948 10548 17000 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17500 10548 17552 10600
rect 17868 10548 17920 10600
rect 18052 10752 18104 10804
rect 18144 10616 18196 10668
rect 16028 10480 16080 10532
rect 18420 10480 18472 10532
rect 15752 10412 15804 10464
rect 17040 10412 17092 10464
rect 17224 10412 17276 10464
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 2504 10208 2556 10260
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 4252 10208 4304 10260
rect 4620 10140 4672 10192
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 2596 10072 2648 10124
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 2504 10004 2556 10056
rect 2688 10004 2740 10056
rect 3792 10004 3844 10056
rect 2228 9979 2280 9988
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2228 9945 2237 9979
rect 2237 9945 2271 9979
rect 2271 9945 2280 9979
rect 2228 9936 2280 9945
rect 4252 9979 4304 9988
rect 4252 9945 4261 9979
rect 4261 9945 4295 9979
rect 4295 9945 4304 9979
rect 5356 10140 5408 10192
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 6368 10208 6420 10260
rect 8024 10251 8076 10260
rect 5632 10072 5684 10124
rect 5080 10004 5132 10013
rect 4252 9936 4304 9945
rect 2596 9868 2648 9920
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3884 9868 3936 9920
rect 4344 9868 4396 9920
rect 4804 9868 4856 9920
rect 5816 9936 5868 9988
rect 6644 10072 6696 10124
rect 7012 10140 7064 10192
rect 7288 10115 7340 10124
rect 6092 10004 6144 10056
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 10968 10208 11020 10260
rect 7840 10140 7892 10192
rect 8208 10140 8260 10192
rect 9312 10140 9364 10192
rect 7472 10004 7524 10056
rect 8392 10072 8444 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9588 10072 9640 10124
rect 8668 10004 8720 10056
rect 6184 9868 6236 9920
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 7196 9868 7248 9920
rect 8208 9936 8260 9988
rect 8300 9936 8352 9988
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 8852 9868 8904 9920
rect 11520 10140 11572 10192
rect 11888 10140 11940 10192
rect 10692 10072 10744 10124
rect 10968 10072 11020 10124
rect 12072 10072 12124 10124
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11888 10004 11940 10056
rect 12532 10140 12584 10192
rect 12808 10115 12860 10124
rect 12808 10081 12817 10115
rect 12817 10081 12851 10115
rect 12851 10081 12860 10115
rect 12808 10072 12860 10081
rect 12992 10072 13044 10124
rect 13360 10004 13412 10056
rect 13544 10004 13596 10056
rect 12624 9979 12676 9988
rect 10508 9911 10560 9920
rect 10508 9877 10517 9911
rect 10517 9877 10551 9911
rect 10551 9877 10560 9911
rect 10508 9868 10560 9877
rect 11244 9868 11296 9920
rect 12624 9945 12633 9979
rect 12633 9945 12667 9979
rect 12667 9945 12676 9979
rect 15752 10140 15804 10192
rect 13912 10072 13964 10124
rect 15108 10072 15160 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 15568 10072 15620 10124
rect 17592 10140 17644 10192
rect 18144 10140 18196 10192
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 15384 10004 15436 10056
rect 12624 9936 12676 9945
rect 13084 9868 13136 9920
rect 15016 9868 15068 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15752 9911 15804 9920
rect 15384 9868 15436 9877
rect 15752 9877 15761 9911
rect 15761 9877 15795 9911
rect 15795 9877 15804 9911
rect 15752 9868 15804 9877
rect 17040 10004 17092 10056
rect 17408 10004 17460 10056
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 17868 10072 17920 10124
rect 18420 10072 18472 10124
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 17960 9936 18012 9988
rect 18512 9936 18564 9988
rect 17776 9868 17828 9920
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 2412 9664 2464 9716
rect 2504 9664 2556 9716
rect 2044 9596 2096 9648
rect 2964 9596 3016 9648
rect 3240 9664 3292 9716
rect 1492 9571 1544 9580
rect 1492 9537 1501 9571
rect 1501 9537 1535 9571
rect 1535 9537 1544 9571
rect 1492 9528 1544 9537
rect 2504 9528 2556 9580
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3148 9528 3200 9580
rect 4436 9596 4488 9648
rect 4804 9664 4856 9716
rect 4988 9596 5040 9648
rect 6000 9664 6052 9716
rect 6368 9664 6420 9716
rect 3976 9528 4028 9580
rect 4252 9528 4304 9580
rect 5908 9596 5960 9648
rect 8300 9664 8352 9716
rect 8944 9664 8996 9716
rect 9312 9707 9364 9716
rect 9312 9673 9321 9707
rect 9321 9673 9355 9707
rect 9355 9673 9364 9707
rect 9312 9664 9364 9673
rect 10232 9664 10284 9716
rect 11244 9664 11296 9716
rect 11980 9707 12032 9716
rect 11980 9673 11989 9707
rect 11989 9673 12023 9707
rect 12023 9673 12032 9707
rect 11980 9664 12032 9673
rect 13084 9664 13136 9716
rect 13360 9664 13412 9716
rect 13912 9664 13964 9716
rect 5816 9528 5868 9580
rect 6644 9528 6696 9580
rect 2044 9460 2096 9512
rect 2228 9392 2280 9444
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 2780 9324 2832 9376
rect 3516 9324 3568 9376
rect 4068 9460 4120 9512
rect 4528 9503 4580 9512
rect 4528 9469 4537 9503
rect 4537 9469 4571 9503
rect 4571 9469 4580 9503
rect 4804 9503 4856 9512
rect 4528 9460 4580 9469
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 6184 9460 6236 9512
rect 6276 9460 6328 9512
rect 4160 9392 4212 9444
rect 4344 9392 4396 9444
rect 4896 9324 4948 9376
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 6000 9392 6052 9444
rect 6368 9435 6420 9444
rect 6368 9401 6377 9435
rect 6377 9401 6411 9435
rect 6411 9401 6420 9435
rect 6368 9392 6420 9401
rect 6828 9460 6880 9512
rect 8024 9528 8076 9580
rect 8576 9596 8628 9648
rect 7196 9460 7248 9512
rect 8300 9460 8352 9512
rect 9128 9528 9180 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 8576 9460 8628 9512
rect 8944 9460 8996 9512
rect 9680 9460 9732 9512
rect 12808 9596 12860 9648
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 10784 9503 10836 9512
rect 8116 9392 8168 9444
rect 8208 9392 8260 9444
rect 9220 9392 9272 9444
rect 10416 9392 10468 9444
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 12440 9528 12492 9580
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 12624 9460 12676 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 13636 9596 13688 9648
rect 14004 9596 14056 9648
rect 14648 9664 14700 9716
rect 15016 9664 15068 9716
rect 15752 9664 15804 9716
rect 16396 9707 16448 9716
rect 16396 9673 16405 9707
rect 16405 9673 16439 9707
rect 16439 9673 16448 9707
rect 16396 9664 16448 9673
rect 16488 9664 16540 9716
rect 18420 9707 18472 9716
rect 14924 9596 14976 9648
rect 15292 9639 15344 9648
rect 15292 9605 15301 9639
rect 15301 9605 15335 9639
rect 15335 9605 15344 9639
rect 15292 9596 15344 9605
rect 15660 9596 15712 9648
rect 17316 9596 17368 9648
rect 17684 9596 17736 9648
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 13084 9460 13136 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 15200 9528 15252 9580
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 15568 9460 15620 9512
rect 16028 9460 16080 9512
rect 18420 9673 18429 9707
rect 18429 9673 18463 9707
rect 18463 9673 18472 9707
rect 18420 9664 18472 9673
rect 17960 9460 18012 9512
rect 6460 9324 6512 9376
rect 6920 9324 6972 9376
rect 10140 9324 10192 9376
rect 10508 9324 10560 9376
rect 11428 9324 11480 9376
rect 11612 9324 11664 9376
rect 13728 9324 13780 9376
rect 14556 9392 14608 9444
rect 17408 9392 17460 9444
rect 17868 9392 17920 9444
rect 18604 9392 18656 9444
rect 14188 9324 14240 9376
rect 14924 9324 14976 9376
rect 18236 9324 18288 9376
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2228 9120 2280 9172
rect 3516 9120 3568 9172
rect 8024 9163 8076 9172
rect 3700 9052 3752 9104
rect 1584 8984 1636 9036
rect 2412 8984 2464 9036
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 4620 9052 4672 9104
rect 4436 9027 4488 9036
rect 1952 8916 2004 8968
rect 1584 8848 1636 8900
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 4712 8984 4764 9036
rect 5632 9027 5684 9036
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 6460 9052 6512 9104
rect 3608 8916 3660 8968
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 8300 9120 8352 9172
rect 9404 9120 9456 9172
rect 9772 9120 9824 9172
rect 9956 9120 10008 9172
rect 11520 9120 11572 9172
rect 14556 9120 14608 9172
rect 9312 9052 9364 9104
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 9496 9027 9548 9036
rect 8668 8984 8720 8993
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 12624 9052 12676 9104
rect 13636 9052 13688 9104
rect 14464 9095 14516 9104
rect 14464 9061 14473 9095
rect 14473 9061 14507 9095
rect 14507 9061 14516 9095
rect 14464 9052 14516 9061
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10048 8984 10100 9036
rect 4896 8848 4948 8900
rect 6828 8891 6880 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2964 8823 3016 8832
rect 2412 8780 2464 8789
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 3240 8780 3292 8832
rect 4068 8780 4120 8832
rect 4436 8780 4488 8832
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5080 8780 5132 8789
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 5908 8780 5960 8832
rect 6828 8857 6862 8891
rect 6862 8857 6880 8891
rect 6828 8848 6880 8857
rect 9772 8916 9824 8968
rect 10140 8916 10192 8968
rect 11244 8984 11296 9036
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11520 9027 11572 9036
rect 11336 8984 11388 8993
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 12440 8984 12492 9036
rect 12808 8984 12860 9036
rect 13544 8984 13596 9036
rect 14556 8984 14608 9036
rect 15200 9120 15252 9172
rect 15292 9120 15344 9172
rect 15752 9120 15804 9172
rect 14924 9052 14976 9104
rect 16948 9052 17000 9104
rect 14832 9027 14884 9036
rect 14832 8993 14841 9027
rect 14841 8993 14875 9027
rect 14875 8993 14884 9027
rect 14832 8984 14884 8993
rect 15016 8984 15068 9036
rect 16120 8984 16172 9036
rect 16304 8984 16356 9036
rect 16856 9027 16908 9036
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 15200 8916 15252 8968
rect 9220 8848 9272 8900
rect 9312 8891 9364 8900
rect 9312 8857 9321 8891
rect 9321 8857 9355 8891
rect 9355 8857 9364 8891
rect 9312 8848 9364 8857
rect 16028 8916 16080 8968
rect 16396 8916 16448 8968
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 16948 8916 17000 8968
rect 7104 8780 7156 8832
rect 8208 8780 8260 8832
rect 9404 8780 9456 8832
rect 9864 8780 9916 8832
rect 11428 8780 11480 8832
rect 12624 8780 12676 8832
rect 14372 8780 14424 8832
rect 14740 8780 14792 8832
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 15384 8780 15436 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 17592 9027 17644 9036
rect 17592 8993 17601 9027
rect 17601 8993 17635 9027
rect 17635 8993 17644 9027
rect 17592 8984 17644 8993
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 17960 8848 18012 8900
rect 18328 8848 18380 8900
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 18512 8780 18564 8832
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 3240 8619 3292 8628
rect 1492 8551 1544 8560
rect 1492 8517 1501 8551
rect 1501 8517 1535 8551
rect 1535 8517 1544 8551
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 3332 8619 3384 8628
rect 3332 8585 3341 8619
rect 3341 8585 3375 8619
rect 3375 8585 3384 8619
rect 4436 8619 4488 8628
rect 3332 8576 3384 8585
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 6828 8576 6880 8628
rect 1492 8508 1544 8517
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 2044 8440 2096 8492
rect 3056 8440 3108 8492
rect 2228 8372 2280 8424
rect 2964 8372 3016 8424
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 2412 8304 2464 8356
rect 4160 8508 4212 8560
rect 3516 8440 3568 8492
rect 4344 8483 4396 8492
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 3884 8304 3936 8356
rect 3516 8236 3568 8288
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 6552 8508 6604 8560
rect 6092 8440 6144 8492
rect 8852 8508 8904 8560
rect 10232 8576 10284 8628
rect 12440 8576 12492 8628
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 13728 8576 13780 8628
rect 15384 8576 15436 8628
rect 15660 8576 15712 8628
rect 16672 8619 16724 8628
rect 16672 8585 16681 8619
rect 16681 8585 16715 8619
rect 16715 8585 16724 8619
rect 16672 8576 16724 8585
rect 17040 8576 17092 8628
rect 17132 8576 17184 8628
rect 17684 8576 17736 8628
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 5908 8372 5960 8424
rect 7472 8483 7524 8492
rect 7472 8449 7506 8483
rect 7506 8449 7524 8483
rect 7472 8440 7524 8449
rect 11152 8508 11204 8560
rect 9220 8440 9272 8492
rect 11336 8440 11388 8492
rect 6644 8372 6696 8424
rect 14832 8440 14884 8492
rect 5816 8304 5868 8356
rect 5908 8236 5960 8288
rect 6184 8236 6236 8288
rect 9036 8304 9088 8356
rect 12716 8304 12768 8356
rect 12992 8347 13044 8356
rect 12992 8313 13001 8347
rect 13001 8313 13035 8347
rect 13035 8313 13044 8347
rect 12992 8304 13044 8313
rect 13176 8347 13228 8356
rect 13176 8313 13185 8347
rect 13185 8313 13219 8347
rect 13219 8313 13228 8347
rect 13176 8304 13228 8313
rect 7932 8236 7984 8288
rect 9404 8236 9456 8288
rect 14464 8372 14516 8424
rect 15292 8508 15344 8560
rect 15568 8508 15620 8560
rect 15476 8440 15528 8492
rect 16764 8440 16816 8492
rect 17500 8440 17552 8492
rect 17960 8440 18012 8492
rect 15936 8304 15988 8356
rect 16396 8304 16448 8356
rect 17500 8304 17552 8356
rect 18880 8372 18932 8424
rect 18788 8304 18840 8356
rect 15108 8236 15160 8288
rect 15660 8236 15712 8288
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 2964 8075 3016 8084
rect 2964 8041 2973 8075
rect 2973 8041 3007 8075
rect 3007 8041 3016 8075
rect 2964 8032 3016 8041
rect 2136 7828 2188 7880
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 3332 7896 3384 7948
rect 4160 7964 4212 8016
rect 4344 8032 4396 8084
rect 5724 8032 5776 8084
rect 5908 8032 5960 8084
rect 3792 7939 3844 7948
rect 3792 7905 3801 7939
rect 3801 7905 3835 7939
rect 3835 7905 3844 7939
rect 3792 7896 3844 7905
rect 4252 7896 4304 7948
rect 4712 7896 4764 7948
rect 4804 7828 4856 7880
rect 5172 7896 5224 7948
rect 7380 8032 7432 8084
rect 7104 7964 7156 8016
rect 9036 7964 9088 8016
rect 15476 8032 15528 8084
rect 15752 8032 15804 8084
rect 17316 8032 17368 8084
rect 17500 8032 17552 8084
rect 18420 8075 18472 8084
rect 18420 8041 18429 8075
rect 18429 8041 18463 8075
rect 18463 8041 18472 8075
rect 18420 8032 18472 8041
rect 14464 7964 14516 8016
rect 5264 7828 5316 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 7564 7896 7616 7948
rect 8852 7828 8904 7880
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 11336 7896 11388 7905
rect 10416 7828 10468 7880
rect 11244 7828 11296 7880
rect 11428 7828 11480 7880
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 15660 7828 15712 7880
rect 17316 7896 17368 7948
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 17592 7896 17644 7905
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 17684 7828 17736 7880
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 18328 7828 18380 7880
rect 3148 7760 3200 7812
rect 3332 7803 3384 7812
rect 3332 7769 3341 7803
rect 3341 7769 3375 7803
rect 3375 7769 3384 7803
rect 3332 7760 3384 7769
rect 4436 7760 4488 7812
rect 5816 7760 5868 7812
rect 7012 7760 7064 7812
rect 10232 7760 10284 7812
rect 10600 7760 10652 7812
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 2044 7692 2096 7744
rect 2504 7692 2556 7744
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 7380 7735 7432 7744
rect 7380 7701 7389 7735
rect 7389 7701 7423 7735
rect 7423 7701 7432 7735
rect 7380 7692 7432 7701
rect 8760 7692 8812 7744
rect 11244 7692 11296 7744
rect 14004 7692 14056 7744
rect 15108 7760 15160 7812
rect 15200 7803 15252 7812
rect 15200 7769 15218 7803
rect 15218 7769 15252 7803
rect 15200 7760 15252 7769
rect 15936 7760 15988 7812
rect 16028 7760 16080 7812
rect 16396 7692 16448 7744
rect 17500 7735 17552 7744
rect 17500 7701 17509 7735
rect 17509 7701 17543 7735
rect 17543 7701 17552 7735
rect 17500 7692 17552 7701
rect 17868 7692 17920 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18236 7692 18288 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 2872 7488 2924 7540
rect 5264 7488 5316 7540
rect 1952 7420 2004 7472
rect 2228 7420 2280 7472
rect 2596 7420 2648 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 2964 7352 3016 7404
rect 3424 7352 3476 7404
rect 2872 7327 2924 7336
rect 1492 7259 1544 7268
rect 1492 7225 1501 7259
rect 1501 7225 1535 7259
rect 1535 7225 1544 7259
rect 1492 7216 1544 7225
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3056 7284 3108 7336
rect 2596 7148 2648 7200
rect 3148 7148 3200 7200
rect 3608 7420 3660 7472
rect 6920 7420 6972 7472
rect 8484 7488 8536 7540
rect 12900 7531 12952 7540
rect 12900 7497 12909 7531
rect 12909 7497 12943 7531
rect 12943 7497 12952 7531
rect 12900 7488 12952 7497
rect 13820 7488 13872 7540
rect 16028 7488 16080 7540
rect 16764 7488 16816 7540
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 8852 7420 8904 7472
rect 4160 7352 4212 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 5540 7395 5592 7404
rect 4344 7352 4396 7361
rect 3700 7284 3752 7336
rect 4068 7216 4120 7268
rect 4712 7284 4764 7336
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 6644 7352 6696 7404
rect 7380 7352 7432 7404
rect 17592 7420 17644 7472
rect 9404 7395 9456 7404
rect 9404 7361 9438 7395
rect 9438 7361 9456 7395
rect 9404 7352 9456 7361
rect 11336 7352 11388 7404
rect 11612 7352 11664 7404
rect 14096 7352 14148 7404
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 15476 7395 15528 7404
rect 5908 7216 5960 7268
rect 12992 7284 13044 7336
rect 13544 7284 13596 7336
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 10692 7216 10744 7268
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16028 7284 16080 7336
rect 17592 7284 17644 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 19064 7284 19116 7336
rect 6828 7148 6880 7200
rect 7564 7148 7616 7200
rect 11244 7148 11296 7200
rect 13452 7148 13504 7200
rect 17408 7216 17460 7268
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 1676 6944 1728 6996
rect 1492 6919 1544 6928
rect 1492 6885 1501 6919
rect 1501 6885 1535 6919
rect 1535 6885 1544 6919
rect 1492 6876 1544 6885
rect 2228 6919 2280 6928
rect 2228 6885 2237 6919
rect 2237 6885 2271 6919
rect 2271 6885 2280 6919
rect 2228 6876 2280 6885
rect 2136 6808 2188 6860
rect 3056 6876 3108 6928
rect 3976 6876 4028 6928
rect 3240 6808 3292 6860
rect 3700 6808 3752 6860
rect 7012 6944 7064 6996
rect 10232 6944 10284 6996
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 1768 6740 1820 6792
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 3056 6740 3108 6792
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 5908 6783 5960 6792
rect 4436 6740 4488 6749
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 3148 6715 3200 6724
rect 3148 6681 3157 6715
rect 3157 6681 3191 6715
rect 3191 6681 3200 6715
rect 3148 6672 3200 6681
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 3332 6604 3384 6656
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4160 6672 4212 6724
rect 4344 6672 4396 6724
rect 5264 6672 5316 6724
rect 5724 6604 5776 6656
rect 6276 6604 6328 6656
rect 7196 6604 7248 6656
rect 8852 6808 8904 6860
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 12992 6851 13044 6860
rect 12992 6817 13001 6851
rect 13001 6817 13035 6851
rect 13035 6817 13044 6851
rect 12992 6808 13044 6817
rect 8668 6740 8720 6792
rect 14832 6944 14884 6996
rect 15108 6944 15160 6996
rect 13728 6876 13780 6928
rect 15936 6944 15988 6996
rect 17316 6944 17368 6996
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 17040 6876 17092 6928
rect 18604 6876 18656 6928
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 17776 6808 17828 6860
rect 18052 6808 18104 6860
rect 8300 6672 8352 6724
rect 9220 6672 9272 6724
rect 11152 6672 11204 6724
rect 11980 6672 12032 6724
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14188 6740 14240 6792
rect 15384 6740 15436 6792
rect 16672 6740 16724 6792
rect 17960 6740 18012 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 8944 6604 8996 6656
rect 10784 6604 10836 6656
rect 12900 6604 12952 6656
rect 13360 6604 13412 6656
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 14832 6672 14884 6724
rect 14280 6604 14332 6656
rect 14648 6604 14700 6656
rect 14740 6604 14792 6656
rect 15936 6672 15988 6724
rect 16120 6672 16172 6724
rect 16212 6604 16264 6656
rect 18328 6672 18380 6724
rect 18420 6604 18472 6656
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 2412 6400 2464 6452
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 3608 6400 3660 6452
rect 2596 6332 2648 6384
rect 4436 6332 4488 6384
rect 12256 6400 12308 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 13176 6400 13228 6452
rect 14096 6400 14148 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 4252 6264 4304 6316
rect 3608 6196 3660 6248
rect 4344 6196 4396 6248
rect 5080 6307 5132 6316
rect 5080 6273 5114 6307
rect 5114 6273 5132 6307
rect 5080 6264 5132 6273
rect 5356 6264 5408 6316
rect 5816 6264 5868 6316
rect 15844 6400 15896 6452
rect 18236 6400 18288 6452
rect 18420 6443 18472 6452
rect 18420 6409 18429 6443
rect 18429 6409 18463 6443
rect 18463 6409 18472 6443
rect 18420 6400 18472 6409
rect 16396 6332 16448 6384
rect 6184 6264 6236 6316
rect 6368 6264 6420 6316
rect 8944 6264 8996 6316
rect 9496 6307 9548 6316
rect 9496 6273 9530 6307
rect 9530 6273 9548 6307
rect 9496 6264 9548 6273
rect 10692 6264 10744 6316
rect 3056 6128 3108 6180
rect 6644 6196 6696 6248
rect 6828 6196 6880 6248
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 10232 6196 10284 6248
rect 11520 6196 11572 6248
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 12808 6264 12860 6316
rect 12900 6264 12952 6316
rect 12992 6196 13044 6248
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 1952 6060 2004 6112
rect 2228 6060 2280 6112
rect 2596 6060 2648 6112
rect 3148 6060 3200 6112
rect 4436 6103 4488 6112
rect 4436 6069 4445 6103
rect 4445 6069 4479 6103
rect 4479 6069 4488 6103
rect 4436 6060 4488 6069
rect 4712 6060 4764 6112
rect 5172 6060 5224 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 6368 6060 6420 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 6736 6103 6788 6112
rect 6736 6069 6745 6103
rect 6745 6069 6779 6103
rect 6779 6069 6788 6103
rect 6736 6060 6788 6069
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 8300 6060 8352 6112
rect 11612 6128 11664 6180
rect 15016 6264 15068 6316
rect 16304 6264 16356 6316
rect 16856 6264 16908 6316
rect 17040 6264 17092 6316
rect 18052 6264 18104 6316
rect 18236 6307 18288 6316
rect 18236 6273 18245 6307
rect 18245 6273 18279 6307
rect 18279 6273 18288 6307
rect 18236 6264 18288 6273
rect 10692 6060 10744 6112
rect 11152 6060 11204 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12624 6060 12676 6112
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 14096 6060 14148 6112
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 17776 6060 17828 6112
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 2872 5856 2924 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4804 5788 4856 5840
rect 1492 5720 1544 5772
rect 2688 5720 2740 5772
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 4528 5720 4580 5772
rect 4620 5720 4672 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 3148 5652 3200 5704
rect 3424 5652 3476 5704
rect 4712 5652 4764 5704
rect 12348 5856 12400 5908
rect 13268 5856 13320 5908
rect 5356 5788 5408 5840
rect 12072 5831 12124 5840
rect 12072 5797 12081 5831
rect 12081 5797 12115 5831
rect 12115 5797 12124 5831
rect 12072 5788 12124 5797
rect 15476 5856 15528 5908
rect 16212 5856 16264 5908
rect 16856 5856 16908 5908
rect 15936 5788 15988 5840
rect 16764 5788 16816 5840
rect 17592 5788 17644 5840
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 11612 5720 11664 5772
rect 12256 5720 12308 5772
rect 6644 5652 6696 5704
rect 6828 5652 6880 5704
rect 8116 5652 8168 5704
rect 9220 5652 9272 5704
rect 1216 5584 1268 5636
rect 3332 5584 3384 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 3700 5516 3752 5568
rect 4436 5516 4488 5568
rect 4620 5516 4672 5568
rect 4988 5516 5040 5568
rect 7104 5584 7156 5636
rect 8208 5516 8260 5568
rect 10232 5652 10284 5704
rect 9312 5584 9364 5636
rect 11336 5652 11388 5704
rect 13912 5652 13964 5704
rect 16396 5720 16448 5772
rect 17408 5720 17460 5772
rect 14188 5652 14240 5704
rect 15108 5652 15160 5704
rect 10692 5584 10744 5636
rect 13084 5584 13136 5636
rect 15200 5584 15252 5636
rect 12348 5516 12400 5568
rect 13728 5516 13780 5568
rect 17316 5652 17368 5704
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 15844 5516 15896 5568
rect 16120 5559 16172 5568
rect 16120 5525 16129 5559
rect 16129 5525 16163 5559
rect 16163 5525 16172 5559
rect 16120 5516 16172 5525
rect 17500 5584 17552 5636
rect 16764 5516 16816 5568
rect 16856 5516 16908 5568
rect 17316 5559 17368 5568
rect 17316 5525 17325 5559
rect 17325 5525 17359 5559
rect 17359 5525 17368 5559
rect 17316 5516 17368 5525
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 3608 5312 3660 5364
rect 3884 5312 3936 5364
rect 4804 5355 4856 5364
rect 4804 5321 4813 5355
rect 4813 5321 4847 5355
rect 4847 5321 4856 5355
rect 4804 5312 4856 5321
rect 9312 5312 9364 5364
rect 9404 5312 9456 5364
rect 1860 5244 1912 5296
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 2228 5176 2280 5228
rect 6276 5244 6328 5296
rect 7380 5244 7432 5296
rect 11980 5312 12032 5364
rect 16304 5312 16356 5364
rect 17316 5312 17368 5364
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 2596 5219 2648 5228
rect 2596 5185 2605 5219
rect 2605 5185 2639 5219
rect 2639 5185 2648 5219
rect 2596 5176 2648 5185
rect 5264 5176 5316 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 7196 5176 7248 5228
rect 8116 5219 8168 5228
rect 2872 5108 2924 5160
rect 3884 5108 3936 5160
rect 4896 5108 4948 5160
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 11336 5244 11388 5296
rect 10232 5219 10284 5228
rect 10232 5185 10266 5219
rect 10266 5185 10284 5219
rect 10232 5176 10284 5185
rect 10692 5176 10744 5228
rect 14188 5244 14240 5296
rect 13728 5176 13780 5228
rect 16948 5244 17000 5296
rect 17500 5244 17552 5296
rect 15660 5176 15712 5228
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 2044 5040 2096 5092
rect 2596 5040 2648 5092
rect 2964 5040 3016 5092
rect 3424 5040 3476 5092
rect 1492 4972 1544 5024
rect 2228 4972 2280 5024
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 3700 4972 3752 5024
rect 4160 5040 4212 5092
rect 4620 5040 4672 5092
rect 5448 5040 5500 5092
rect 6276 4972 6328 5024
rect 8760 4972 8812 5024
rect 9588 4972 9640 5024
rect 16580 5176 16632 5228
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 17316 5108 17368 5160
rect 18604 5176 18656 5228
rect 18972 5108 19024 5160
rect 11428 4972 11480 5024
rect 11980 4972 12032 5024
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 18328 5040 18380 5092
rect 18236 4972 18288 5024
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3884 4768 3936 4820
rect 4528 4768 4580 4820
rect 4804 4768 4856 4820
rect 6092 4768 6144 4820
rect 6828 4768 6880 4820
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 2780 4632 2832 4684
rect 3424 4700 3476 4752
rect 4068 4700 4120 4752
rect 8024 4768 8076 4820
rect 11428 4768 11480 4820
rect 14740 4768 14792 4820
rect 15200 4768 15252 4820
rect 13728 4700 13780 4752
rect 2596 4564 2648 4616
rect 3056 4564 3108 4616
rect 4160 4564 4212 4616
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 5080 4564 5132 4616
rect 5448 4607 5500 4616
rect 5448 4573 5466 4607
rect 5466 4573 5500 4607
rect 5448 4564 5500 4573
rect 6644 4564 6696 4616
rect 10140 4607 10192 4616
rect 10140 4573 10158 4607
rect 10158 4573 10192 4607
rect 10600 4607 10652 4616
rect 10140 4564 10192 4573
rect 3148 4496 3200 4548
rect 6368 4496 6420 4548
rect 7012 4496 7064 4548
rect 7288 4496 7340 4548
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2412 4471 2464 4480
rect 2412 4437 2421 4471
rect 2421 4437 2455 4471
rect 2455 4437 2464 4471
rect 2412 4428 2464 4437
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 3884 4428 3936 4480
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 4712 4428 4764 4480
rect 5172 4428 5224 4480
rect 7472 4428 7524 4480
rect 9588 4496 9640 4548
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 11796 4564 11848 4616
rect 16764 4768 16816 4820
rect 17040 4768 17092 4820
rect 18144 4768 18196 4820
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 15568 4700 15620 4752
rect 16396 4700 16448 4752
rect 16856 4632 16908 4684
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 11520 4496 11572 4548
rect 12256 4496 12308 4548
rect 15752 4564 15804 4616
rect 17132 4564 17184 4616
rect 17868 4632 17920 4684
rect 19064 4632 19116 4684
rect 17684 4564 17736 4616
rect 18052 4564 18104 4616
rect 12440 4428 12492 4480
rect 13084 4471 13136 4480
rect 13084 4437 13093 4471
rect 13093 4437 13127 4471
rect 13127 4437 13136 4471
rect 13084 4428 13136 4437
rect 15108 4496 15160 4548
rect 16028 4496 16080 4548
rect 17408 4496 17460 4548
rect 15936 4428 15988 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 16396 4471 16448 4480
rect 16396 4437 16405 4471
rect 16405 4437 16439 4471
rect 16439 4437 16448 4471
rect 16396 4428 16448 4437
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 1308 4224 1360 4276
rect 2596 4224 2648 4276
rect 3056 4224 3108 4276
rect 5724 4224 5776 4276
rect 11796 4267 11848 4276
rect 3424 4199 3476 4208
rect 1860 4088 1912 4140
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 3424 4165 3433 4199
rect 3433 4165 3467 4199
rect 3467 4165 3476 4199
rect 3424 4156 3476 4165
rect 4528 4156 4580 4208
rect 8024 4156 8076 4208
rect 3056 4131 3108 4140
rect 1492 3995 1544 4004
rect 1492 3961 1501 3995
rect 1501 3961 1535 3995
rect 1535 3961 1544 3995
rect 1492 3952 1544 3961
rect 2044 3952 2096 4004
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 2504 4020 2556 4072
rect 4712 4088 4764 4140
rect 5080 4131 5132 4140
rect 5080 4097 5114 4131
rect 5114 4097 5132 4131
rect 5080 4088 5132 4097
rect 5908 4088 5960 4140
rect 6552 4088 6604 4140
rect 8208 4088 8260 4140
rect 8392 4088 8444 4140
rect 11796 4233 11805 4267
rect 11805 4233 11839 4267
rect 11839 4233 11848 4267
rect 11796 4224 11848 4233
rect 12256 4224 12308 4276
rect 13084 4224 13136 4276
rect 15568 4224 15620 4276
rect 16396 4224 16448 4276
rect 16948 4224 17000 4276
rect 18512 4224 18564 4276
rect 11336 4156 11388 4208
rect 11244 4088 11296 4140
rect 11428 4088 11480 4140
rect 11704 4088 11756 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12716 4131 12768 4140
rect 12716 4097 12750 4131
rect 12750 4097 12768 4131
rect 3148 3952 3200 4004
rect 4712 3952 4764 4004
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 1952 3884 2004 3936
rect 2320 3884 2372 3936
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 4252 3884 4304 3936
rect 7012 3952 7064 4004
rect 8116 3952 8168 4004
rect 5724 3884 5776 3936
rect 6276 3884 6328 3936
rect 8760 3884 8812 3936
rect 11612 3952 11664 4004
rect 12716 4088 12768 4097
rect 13544 4088 13596 4140
rect 15200 4156 15252 4208
rect 16120 4156 16172 4208
rect 16764 4156 16816 4208
rect 13820 4020 13872 4072
rect 17224 4088 17276 4140
rect 17592 4199 17644 4208
rect 17592 4165 17601 4199
rect 17601 4165 17635 4199
rect 17635 4165 17644 4199
rect 17592 4156 17644 4165
rect 15292 4020 15344 4072
rect 15660 4063 15712 4072
rect 15660 4029 15669 4063
rect 15669 4029 15703 4063
rect 15703 4029 15712 4063
rect 15660 4020 15712 4029
rect 16212 4020 16264 4072
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 12348 3927 12400 3936
rect 12348 3893 12357 3927
rect 12357 3893 12391 3927
rect 12391 3893 12400 3927
rect 12348 3884 12400 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 17316 4020 17368 4072
rect 18696 4088 18748 4140
rect 18880 4020 18932 4072
rect 17040 3952 17092 4004
rect 17960 3995 18012 4004
rect 17960 3961 17969 3995
rect 17969 3961 18003 3995
rect 18003 3961 18012 3995
rect 17960 3952 18012 3961
rect 15292 3884 15344 3936
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 4160 3680 4212 3732
rect 4712 3680 4764 3732
rect 8576 3680 8628 3732
rect 6552 3655 6604 3664
rect 1952 3544 2004 3596
rect 3056 3587 3108 3596
rect 3056 3553 3065 3587
rect 3065 3553 3099 3587
rect 3099 3553 3108 3587
rect 3056 3544 3108 3553
rect 3332 3544 3384 3596
rect 4436 3544 4488 3596
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 2228 3476 2280 3528
rect 2688 3476 2740 3528
rect 2780 3476 2832 3528
rect 3516 3476 3568 3528
rect 4344 3476 4396 3528
rect 6552 3621 6561 3655
rect 6561 3621 6595 3655
rect 6595 3621 6604 3655
rect 6552 3612 6604 3621
rect 8208 3544 8260 3596
rect 5724 3476 5776 3528
rect 6184 3476 6236 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 2228 3340 2280 3392
rect 2412 3340 2464 3392
rect 4712 3408 4764 3460
rect 4896 3408 4948 3460
rect 8116 3408 8168 3460
rect 8484 3476 8536 3528
rect 11060 3680 11112 3732
rect 10324 3612 10376 3664
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 9772 3476 9824 3528
rect 15200 3680 15252 3732
rect 12348 3612 12400 3664
rect 12532 3544 12584 3596
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 15752 3680 15804 3732
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 17408 3680 17460 3732
rect 18328 3723 18380 3732
rect 18328 3689 18337 3723
rect 18337 3689 18371 3723
rect 18371 3689 18380 3723
rect 18328 3680 18380 3689
rect 17776 3612 17828 3664
rect 17684 3544 17736 3596
rect 4344 3383 4396 3392
rect 4344 3349 4353 3383
rect 4353 3349 4387 3383
rect 4387 3349 4396 3383
rect 4344 3340 4396 3349
rect 4528 3340 4580 3392
rect 5172 3340 5224 3392
rect 7932 3340 7984 3392
rect 8024 3340 8076 3392
rect 8392 3340 8444 3392
rect 8760 3340 8812 3392
rect 9312 3408 9364 3460
rect 11980 3476 12032 3528
rect 12900 3476 12952 3528
rect 12992 3476 13044 3528
rect 16212 3476 16264 3528
rect 18788 3544 18840 3596
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 10876 3340 10928 3392
rect 11796 3340 11848 3392
rect 12348 3408 12400 3460
rect 13084 3408 13136 3460
rect 13452 3408 13504 3460
rect 12716 3340 12768 3392
rect 12808 3340 12860 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 15384 3408 15436 3460
rect 15568 3408 15620 3460
rect 17960 3408 18012 3460
rect 18972 3476 19024 3528
rect 17776 3340 17828 3392
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 4252 3179 4304 3188
rect 2780 3068 2832 3120
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 4620 3136 4672 3188
rect 5080 3136 5132 3188
rect 9312 3136 9364 3188
rect 9772 3136 9824 3188
rect 1676 3000 1728 3052
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 3332 3000 3384 3052
rect 3424 3043 3476 3052
rect 3424 3009 3433 3043
rect 3433 3009 3467 3043
rect 3467 3009 3476 3043
rect 3700 3043 3752 3052
rect 3424 3000 3476 3009
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 5816 3068 5868 3120
rect 6184 3068 6236 3120
rect 3884 2932 3936 2984
rect 2964 2864 3016 2916
rect 1400 2839 1452 2848
rect 1400 2805 1409 2839
rect 1409 2805 1443 2839
rect 1443 2805 1452 2839
rect 1400 2796 1452 2805
rect 1676 2796 1728 2848
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 2780 2796 2832 2848
rect 3976 2864 4028 2916
rect 4620 2932 4672 2984
rect 4804 3000 4856 3052
rect 6092 3000 6144 3052
rect 7104 3000 7156 3052
rect 8208 3068 8260 3120
rect 5172 2932 5224 2984
rect 6184 2975 6236 2984
rect 6184 2941 6193 2975
rect 6193 2941 6227 2975
rect 6227 2941 6236 2975
rect 6184 2932 6236 2941
rect 4988 2864 5040 2916
rect 8116 2932 8168 2984
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 8576 3000 8628 3052
rect 11336 3068 11388 3120
rect 10048 3000 10100 3052
rect 10232 3043 10284 3052
rect 10232 3009 10266 3043
rect 10266 3009 10284 3043
rect 10232 3000 10284 3009
rect 11796 3136 11848 3188
rect 12440 3136 12492 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13728 3068 13780 3120
rect 13820 3068 13872 3120
rect 13268 3000 13320 3052
rect 13544 3000 13596 3052
rect 15476 3068 15528 3120
rect 16028 3136 16080 3188
rect 16856 3136 16908 3188
rect 17132 3136 17184 3188
rect 18512 3136 18564 3188
rect 15568 3000 15620 3052
rect 16396 3000 16448 3052
rect 17592 3000 17644 3052
rect 8300 2932 8352 2984
rect 3608 2839 3660 2848
rect 3608 2805 3617 2839
rect 3617 2805 3651 2839
rect 3651 2805 3660 2839
rect 4712 2839 4764 2848
rect 3608 2796 3660 2805
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 7196 2796 7248 2848
rect 8116 2796 8168 2848
rect 8668 2796 8720 2848
rect 9220 2796 9272 2848
rect 9680 2796 9732 2848
rect 10324 2796 10376 2848
rect 11152 2864 11204 2916
rect 17776 2932 17828 2984
rect 11428 2796 11480 2848
rect 17960 2864 18012 2916
rect 13176 2796 13228 2848
rect 13636 2796 13688 2848
rect 15568 2796 15620 2848
rect 16856 2796 16908 2848
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 3884 2635 3936 2644
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 5264 2592 5316 2644
rect 9128 2635 9180 2644
rect 1216 2524 1268 2576
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 2320 2388 2372 2440
rect 2872 2456 2924 2508
rect 3700 2524 3752 2576
rect 4712 2524 4764 2576
rect 4068 2456 4120 2508
rect 2964 2320 3016 2372
rect 3608 2388 3660 2440
rect 4988 2456 5040 2508
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 9588 2592 9640 2644
rect 11520 2635 11572 2644
rect 9496 2524 9548 2576
rect 11520 2601 11529 2635
rect 11529 2601 11563 2635
rect 11563 2601 11572 2635
rect 11520 2592 11572 2601
rect 11980 2592 12032 2644
rect 14740 2592 14792 2644
rect 16212 2592 16264 2644
rect 17776 2592 17828 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 18420 2635 18472 2644
rect 18420 2601 18429 2635
rect 18429 2601 18463 2635
rect 18463 2601 18472 2635
rect 18420 2592 18472 2601
rect 13176 2567 13228 2576
rect 13176 2533 13185 2567
rect 13185 2533 13219 2567
rect 13219 2533 13228 2567
rect 13176 2524 13228 2533
rect 15568 2524 15620 2576
rect 4804 2388 4856 2440
rect 6000 2431 6052 2440
rect 4620 2320 4672 2372
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 1860 2252 1912 2261
rect 2044 2252 2096 2304
rect 2872 2252 2924 2304
rect 3700 2252 3752 2304
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 6460 2388 6512 2440
rect 11336 2499 11388 2508
rect 8300 2388 8352 2440
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 10048 2388 10100 2440
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 13268 2456 13320 2508
rect 12992 2431 13044 2440
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 6920 2252 6972 2304
rect 7288 2320 7340 2372
rect 7380 2320 7432 2372
rect 9220 2320 9272 2372
rect 9404 2320 9456 2372
rect 7932 2252 7984 2304
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 13084 2388 13136 2440
rect 9772 2252 9824 2304
rect 10692 2252 10744 2304
rect 14096 2456 14148 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 16856 2456 16908 2508
rect 16304 2388 16356 2440
rect 17408 2431 17460 2440
rect 14648 2320 14700 2372
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 14832 2252 14884 2304
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17868 2431 17920 2440
rect 17500 2388 17552 2397
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 18144 2388 18196 2440
rect 16948 2295 17000 2304
rect 16948 2261 16957 2295
rect 16957 2261 16991 2295
rect 16991 2261 17000 2295
rect 16948 2252 17000 2261
rect 17776 2252 17828 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 1492 2048 1544 2100
rect 4620 2048 4672 2100
rect 7380 2048 7432 2100
rect 14188 2048 14240 2100
rect 17868 2048 17920 2100
rect 6552 1980 6604 2032
rect 12992 1980 13044 2032
rect 13360 1980 13412 2032
rect 16948 1980 17000 2032
rect 3056 1912 3108 1964
rect 7932 1912 7984 1964
rect 8116 1912 8168 1964
rect 14096 1912 14148 1964
rect 9772 1844 9824 1896
rect 12716 1776 12768 1828
rect 15384 1776 15436 1828
<< metal2 >>
rect 1122 16400 1178 17200
rect 3330 16400 3386 17200
rect 4434 16688 4490 16697
rect 4434 16623 4490 16632
rect 1136 13802 1164 16400
rect 2962 15464 3018 15473
rect 2962 15399 3018 15408
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1124 13796 1176 13802
rect 1124 13738 1176 13744
rect 1216 13184 1268 13190
rect 1216 13126 1268 13132
rect 1124 11552 1176 11558
rect 1124 11494 1176 11500
rect 1136 3369 1164 11494
rect 1228 5642 1256 13126
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1504 11393 1532 11698
rect 1490 11384 1546 11393
rect 1490 11319 1546 11328
rect 1490 10568 1546 10577
rect 1490 10503 1546 10512
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1306 8392 1362 8401
rect 1306 8327 1362 8336
rect 1216 5636 1268 5642
rect 1216 5578 1268 5584
rect 1320 4282 1348 8327
rect 1412 5710 1440 10406
rect 1504 10062 1532 10503
rect 1492 10056 1544 10062
rect 1688 10033 1716 11698
rect 1780 11354 1808 13806
rect 1964 12345 1992 14350
rect 2240 14249 2268 14418
rect 2226 14240 2282 14249
rect 2226 14175 2282 14184
rect 2226 13832 2282 13841
rect 2332 13818 2360 14962
rect 2778 14648 2834 14657
rect 2778 14583 2780 14592
rect 2832 14583 2834 14592
rect 2780 14554 2832 14560
rect 2792 14482 2820 14554
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2976 14414 3004 15399
rect 3054 15056 3110 15065
rect 3054 14991 3110 15000
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 13938 3004 14350
rect 3068 14346 3096 14991
rect 3344 14906 3372 16400
rect 3698 16280 3754 16289
rect 3698 16215 3754 16224
rect 3606 15872 3662 15881
rect 3606 15807 3662 15816
rect 3344 14878 3556 14906
rect 3620 14890 3648 15807
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 3528 14482 3556 14878
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2282 13790 2360 13818
rect 2226 13767 2282 13776
rect 2240 13326 2268 13767
rect 2792 13433 2820 13874
rect 2872 13864 2924 13870
rect 2870 13832 2872 13841
rect 2924 13832 2926 13841
rect 3160 13818 3188 14214
rect 3344 13977 3372 14214
rect 3620 14056 3648 14826
rect 3436 14028 3648 14056
rect 3330 13968 3386 13977
rect 3330 13903 3386 13912
rect 3436 13870 3464 14028
rect 3712 13954 3740 16215
rect 4448 14822 4476 16623
rect 5538 16538 5594 17200
rect 7746 16538 7802 17200
rect 5538 16510 5764 16538
rect 5538 16400 5594 16510
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 4448 14414 4476 14758
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4894 14376 4950 14385
rect 3528 13938 3740 13954
rect 4080 13938 4108 14350
rect 3528 13932 3752 13938
rect 3528 13926 3700 13932
rect 2870 13767 2926 13776
rect 2976 13790 3188 13818
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 2778 13424 2834 13433
rect 2778 13359 2834 13368
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 1950 12336 2006 12345
rect 1950 12271 2006 12280
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1492 9998 1544 10004
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 1584 9920 1636 9926
rect 1490 9888 1546 9897
rect 1584 9862 1636 9868
rect 1490 9823 1546 9832
rect 1504 9586 1532 9823
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1596 9042 1624 9862
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1584 8900 1636 8906
rect 1504 8566 1532 8871
rect 1584 8842 1636 8848
rect 1596 8634 1624 8842
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1492 8560 1544 8566
rect 1688 8514 1716 9959
rect 1768 8832 1820 8838
rect 1766 8800 1768 8809
rect 1820 8800 1822 8809
rect 1766 8735 1822 8744
rect 1766 8664 1822 8673
rect 1766 8599 1822 8608
rect 1492 8502 1544 8508
rect 1596 8486 1716 8514
rect 1780 8498 1808 8599
rect 1768 8492 1820 8498
rect 1490 8120 1546 8129
rect 1490 8055 1492 8064
rect 1544 8055 1546 8064
rect 1492 8026 1544 8032
rect 1490 7304 1546 7313
rect 1490 7239 1492 7248
rect 1544 7239 1546 7248
rect 1492 7210 1544 7216
rect 1492 6928 1544 6934
rect 1490 6896 1492 6905
rect 1544 6896 1546 6905
rect 1490 6831 1546 6840
rect 1596 6202 1624 8486
rect 1768 8434 1820 8440
rect 1872 7834 1900 11222
rect 1964 11121 1992 12174
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 2056 11801 2084 12106
rect 2042 11792 2098 11801
rect 2042 11727 2098 11736
rect 2148 11744 2176 12922
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2240 12617 2268 12718
rect 2226 12608 2282 12617
rect 2226 12543 2282 12552
rect 2228 12232 2280 12238
rect 2226 12200 2228 12209
rect 2280 12200 2282 12209
rect 2226 12135 2282 12144
rect 2148 11716 2360 11744
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1950 11112 2006 11121
rect 1950 11047 2006 11056
rect 1964 10810 1992 11047
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9178 1992 10542
rect 2056 9654 2084 11630
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 8362 1992 8910
rect 2056 8634 2084 9454
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 2056 7993 2084 8434
rect 2042 7984 2098 7993
rect 2042 7919 2098 7928
rect 2148 7886 2176 11562
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10985 2268 11086
rect 2226 10976 2282 10985
rect 2226 10911 2282 10920
rect 2240 10742 2268 10911
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2332 10674 2360 11716
rect 2424 11218 2452 12718
rect 2516 11626 2544 12786
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2608 11898 2636 12718
rect 2700 12238 2728 13126
rect 2884 13025 2912 13194
rect 2976 13190 3004 13790
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 3068 13530 3096 13670
rect 3174 13628 3482 13637
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13563 3482 13572
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2870 13016 2926 13025
rect 2870 12951 2926 12960
rect 2976 12889 3004 13126
rect 3068 12986 3096 13330
rect 3436 13326 3464 13466
rect 3148 13320 3200 13326
rect 3146 13288 3148 13297
rect 3424 13320 3476 13326
rect 3200 13288 3202 13297
rect 3424 13262 3476 13268
rect 3146 13223 3202 13232
rect 3528 12986 3556 13926
rect 3700 13874 3752 13880
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3974 13832 4030 13841
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 2962 12880 3018 12889
rect 2962 12815 3018 12824
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2792 12102 2820 12650
rect 2976 12481 3004 12650
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 2962 12472 3018 12481
rect 3174 12475 3482 12484
rect 2872 12436 2924 12442
rect 2962 12407 3018 12416
rect 2872 12378 2924 12384
rect 2884 12186 2912 12378
rect 3528 12306 3556 12582
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3528 12209 3556 12242
rect 3514 12200 3570 12209
rect 2884 12158 3004 12186
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2792 11801 2820 12038
rect 2778 11792 2834 11801
rect 2778 11727 2834 11736
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2502 11248 2558 11257
rect 2412 11212 2464 11218
rect 2502 11183 2558 11192
rect 2412 11154 2464 11160
rect 2424 10985 2452 11154
rect 2516 11150 2544 11183
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2410 10976 2466 10985
rect 2410 10911 2466 10920
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2240 9761 2268 9930
rect 2226 9752 2282 9761
rect 2226 9687 2282 9696
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2240 9178 2268 9386
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2332 8786 2360 10610
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 9722 2452 10406
rect 2516 10266 2544 11086
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2700 10810 2728 11018
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2516 9722 2544 9998
rect 2608 9926 2636 10066
rect 2700 10062 2728 10610
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2504 9716 2556 9722
rect 2792 9674 2820 11630
rect 2884 9761 2912 12038
rect 2870 9752 2926 9761
rect 2976 9738 3004 12158
rect 3514 12135 3570 12144
rect 3054 11792 3110 11801
rect 3054 11727 3110 11736
rect 3068 11150 3096 11727
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 11558 3556 11630
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3068 10713 3096 10746
rect 3054 10704 3110 10713
rect 3160 10674 3188 10950
rect 3054 10639 3110 10648
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3528 10606 3556 11494
rect 3620 10713 3648 13806
rect 3804 13569 3832 13806
rect 3974 13767 4030 13776
rect 4068 13796 4120 13802
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3790 13560 3846 13569
rect 3790 13495 3846 13504
rect 3698 13424 3754 13433
rect 3896 13394 3924 13670
rect 3698 13359 3754 13368
rect 3884 13388 3936 13394
rect 3712 13258 3740 13359
rect 3884 13330 3936 13336
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3896 12986 3924 13330
rect 3988 13190 4016 13767
rect 4068 13738 4120 13744
rect 4080 13433 4108 13738
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 4158 13288 4214 13297
rect 4158 13223 4160 13232
rect 4212 13223 4214 13232
rect 4160 13194 4212 13200
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3606 10704 3662 10713
rect 3606 10639 3662 10648
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 10266 3096 10474
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3068 10169 3096 10202
rect 3054 10160 3110 10169
rect 3054 10095 3110 10104
rect 3148 9920 3200 9926
rect 3528 9897 3556 10542
rect 3606 10432 3662 10441
rect 3606 10367 3662 10376
rect 3148 9862 3200 9868
rect 3514 9888 3570 9897
rect 2976 9710 3096 9738
rect 2870 9687 2926 9696
rect 2504 9658 2556 9664
rect 2700 9646 2820 9674
rect 2964 9648 3016 9654
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 8945 2452 8978
rect 2410 8936 2466 8945
rect 2410 8871 2466 8880
rect 2424 8838 2452 8871
rect 2240 8758 2360 8786
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2240 8430 2268 8758
rect 2318 8664 2374 8673
rect 2318 8599 2374 8608
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2332 7886 2360 8599
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 1780 7806 1900 7834
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1688 7002 1716 7346
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1780 6882 1808 7806
rect 1860 7744 1912 7750
rect 1858 7712 1860 7721
rect 2044 7744 2096 7750
rect 1912 7712 1914 7721
rect 2044 7686 2096 7692
rect 1858 7647 1914 7656
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1688 6854 1808 6882
rect 1688 6322 1716 6854
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1780 6458 1808 6734
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6497 1900 6598
rect 1858 6488 1914 6497
rect 1768 6452 1820 6458
rect 1858 6423 1914 6432
rect 1768 6394 1820 6400
rect 1964 6322 1992 7414
rect 2056 6798 2084 7686
rect 2228 7472 2280 7478
rect 2226 7440 2228 7449
rect 2280 7440 2282 7449
rect 2136 7404 2188 7410
rect 2226 7375 2282 7384
rect 2136 7346 2188 7352
rect 2148 6866 2176 7346
rect 2332 7324 2360 7822
rect 2240 7296 2360 7324
rect 2240 6934 2268 7296
rect 2228 6928 2280 6934
rect 2228 6870 2280 6876
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2424 6458 2452 8298
rect 2516 7750 2544 9522
rect 2700 9382 2728 9646
rect 3068 9625 3096 9710
rect 2964 9590 3016 9596
rect 3054 9616 3110 9625
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2780 9376 2832 9382
rect 2884 9353 2912 9522
rect 2976 9466 3004 9590
rect 3160 9586 3188 9862
rect 3514 9823 3570 9832
rect 3240 9716 3292 9722
rect 3620 9674 3648 10367
rect 3240 9658 3292 9664
rect 3054 9551 3110 9560
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3252 9466 3280 9658
rect 2976 9438 3280 9466
rect 3528 9646 3648 9674
rect 3712 9674 3740 12242
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3790 11384 3846 11393
rect 3790 11319 3792 11328
rect 3844 11319 3846 11328
rect 3792 11290 3844 11296
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9738 3832 9998
rect 3896 9926 3924 11834
rect 3988 11082 4016 12650
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12238 4200 12582
rect 4264 12442 4292 14350
rect 4894 14311 4950 14320
rect 4908 14278 4936 14311
rect 5460 14278 5488 14758
rect 5736 14618 5764 16510
rect 7484 16510 7802 16538
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5552 14414 5580 14486
rect 5920 14414 5948 14894
rect 6564 14618 6592 14962
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4342 12744 4398 12753
rect 4342 12679 4398 12688
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4068 12096 4120 12102
rect 4356 12050 4384 12679
rect 4068 12038 4120 12044
rect 4080 11898 4108 12038
rect 4172 12022 4384 12050
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4172 11762 4200 12022
rect 4448 11880 4476 14010
rect 5000 13870 5028 14214
rect 5276 14074 5304 14214
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 6932 14074 6960 14826
rect 7484 14618 7512 16510
rect 7746 16400 7802 16510
rect 9954 16538 10010 17200
rect 12162 16538 12218 17200
rect 9954 16510 10180 16538
rect 9954 16400 10010 16510
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 10152 14618 10180 16510
rect 11992 16510 12218 16538
rect 11992 14618 12020 16510
rect 12162 16400 12218 16510
rect 14370 16538 14426 17200
rect 16302 16552 16358 16561
rect 14370 16510 14596 16538
rect 14370 16400 14426 16510
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 14568 14618 14596 16510
rect 16302 16487 16358 16496
rect 16578 16538 16634 17200
rect 16578 16510 16896 16538
rect 16026 16144 16082 16153
rect 16026 16079 16082 16088
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 15212 14482 15240 14758
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6012 13870 6040 14010
rect 7378 13968 7434 13977
rect 7378 13903 7434 13912
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 4632 13530 4660 13806
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4724 13410 4752 13806
rect 4896 13728 4948 13734
rect 5092 13682 5120 13806
rect 6460 13728 6512 13734
rect 4948 13676 5120 13682
rect 4896 13670 5120 13676
rect 4908 13654 5120 13670
rect 5722 13696 5778 13705
rect 6460 13670 6512 13676
rect 5722 13631 5778 13640
rect 4632 13382 4752 13410
rect 4894 13424 4950 13433
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12986 4568 13126
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4540 12306 4568 12718
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4356 11852 4476 11880
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4356 11676 4384 11852
rect 4528 11688 4580 11694
rect 4356 11648 4476 11676
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3974 10840 4030 10849
rect 3974 10775 3976 10784
rect 4028 10775 4030 10784
rect 3976 10746 4028 10752
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3974 9752 4030 9761
rect 3804 9710 3974 9738
rect 3974 9687 4030 9696
rect 3712 9646 3924 9674
rect 2780 9318 2832 9324
rect 2870 9344 2926 9353
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2608 7478 2636 8978
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2502 6896 2558 6905
rect 2502 6831 2558 6840
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2516 6322 2544 6831
rect 2608 6390 2636 7142
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2240 6225 2268 6258
rect 2226 6216 2282 6225
rect 1596 6174 1900 6202
rect 1492 6112 1544 6118
rect 1490 6080 1492 6089
rect 1544 6080 1546 6089
rect 1490 6015 1546 6024
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1504 5522 1532 5714
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1596 5574 1624 5607
rect 1412 5494 1532 5522
rect 1584 5568 1636 5574
rect 1768 5568 1820 5574
rect 1584 5510 1636 5516
rect 1674 5536 1730 5545
rect 1308 4276 1360 4282
rect 1308 4218 1360 4224
rect 1122 3360 1178 3369
rect 1122 3295 1178 3304
rect 1412 3074 1440 5494
rect 1768 5510 1820 5516
rect 1674 5471 1730 5480
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1504 5273 1532 5306
rect 1490 5264 1546 5273
rect 1688 5234 1716 5471
rect 1490 5199 1546 5208
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4865 1532 4966
rect 1490 4856 1546 4865
rect 1490 4791 1546 4800
rect 1492 4480 1544 4486
rect 1490 4448 1492 4457
rect 1544 4448 1546 4457
rect 1490 4383 1546 4392
rect 1490 4040 1546 4049
rect 1490 3975 1492 3984
rect 1544 3975 1546 3984
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1492 3946 1544 3952
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 3233 1532 3334
rect 1490 3224 1546 3233
rect 1490 3159 1546 3168
rect 1412 3046 1532 3074
rect 1688 3058 1716 3975
rect 1780 3534 1808 5510
rect 1872 5302 1900 6174
rect 2226 6151 2282 6160
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 1964 4808 1992 6054
rect 2134 5264 2190 5273
rect 2240 5234 2268 6054
rect 2134 5199 2190 5208
rect 2228 5228 2280 5234
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1872 4780 1992 4808
rect 1872 4146 1900 4780
rect 1950 4720 2006 4729
rect 1950 4655 2006 4664
rect 1964 4622 1992 4655
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 2056 4146 2084 5034
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1952 3936 2004 3942
rect 2056 3913 2084 3946
rect 1952 3878 2004 3884
rect 2042 3904 2098 3913
rect 1872 3641 1900 3878
rect 1858 3632 1914 3641
rect 1964 3602 1992 3878
rect 2042 3839 2098 3848
rect 1858 3567 1914 3576
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1216 2576 1268 2582
rect 1216 2518 1268 2524
rect 1228 800 1256 2518
rect 1412 2446 1440 2790
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1504 2106 1532 3046
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1676 2848 1728 2854
rect 1582 2816 1638 2825
rect 1676 2790 1728 2796
rect 1582 2751 1638 2760
rect 1596 2650 1624 2751
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1492 2100 1544 2106
rect 1492 2042 1544 2048
rect 1214 0 1270 800
rect 1688 785 1716 2790
rect 1858 2408 1914 2417
rect 1858 2343 1914 2352
rect 1872 2310 1900 2343
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1964 1193 1992 3334
rect 2056 2825 2084 3839
rect 2148 3058 2176 5199
rect 2228 5170 2280 5176
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2240 3534 2268 4966
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2042 2816 2098 2825
rect 2042 2751 2098 2760
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1950 1184 2006 1193
rect 1950 1119 2006 1128
rect 2056 800 2084 2246
rect 2240 2009 2268 3334
rect 2332 2446 2360 3878
rect 2424 3398 2452 4422
rect 2516 4078 2544 6258
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5234 2636 6054
rect 2700 5778 2728 9318
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2792 5624 2820 9318
rect 2870 9279 2926 9288
rect 2976 9194 3004 9438
rect 3528 9382 3556 9646
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 2884 9166 3004 9194
rect 3528 9178 3556 9318
rect 3516 9172 3568 9178
rect 2884 7546 2912 9166
rect 3516 9114 3568 9120
rect 3330 9072 3386 9081
rect 3330 9007 3386 9016
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 2976 8537 3004 8774
rect 3252 8634 3280 8774
rect 3344 8634 3372 9007
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 2962 8528 3018 8537
rect 3528 8498 3556 9114
rect 3620 8974 3648 9415
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 2962 8463 3018 8472
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 8090 3004 8366
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2884 5914 2912 7278
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2700 5596 2820 5624
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2608 5098 2636 5170
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2608 4282 2636 4558
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2608 3505 2636 4218
rect 2700 3534 2728 5596
rect 2976 5250 3004 7346
rect 3068 7342 3096 8434
rect 3424 8424 3476 8430
rect 3422 8392 3424 8401
rect 3476 8392 3478 8401
rect 3422 8327 3478 8336
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7818 3372 7890
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3056 7336 3108 7342
rect 3160 7313 3188 7754
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7410 3464 7686
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3056 7278 3108 7284
rect 3146 7304 3202 7313
rect 3146 7239 3202 7248
rect 3148 7200 3200 7206
rect 3068 7160 3148 7188
rect 3068 6934 3096 7160
rect 3148 7142 3200 7148
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6186 3096 6734
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3160 6118 3188 6666
rect 3252 6458 3280 6802
rect 3330 6760 3386 6769
rect 3330 6695 3386 6704
rect 3344 6662 3372 6695
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 3146 5808 3202 5817
rect 3056 5772 3108 5778
rect 3146 5743 3202 5752
rect 3056 5714 3108 5720
rect 3068 5681 3096 5714
rect 3160 5710 3188 5743
rect 3148 5704 3200 5710
rect 3054 5672 3110 5681
rect 3148 5646 3200 5652
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3054 5607 3110 5616
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 2976 5222 3096 5250
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4690 2820 4966
rect 2884 4826 2912 5102
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 3534 2820 4422
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2688 3528 2740 3534
rect 2594 3496 2650 3505
rect 2688 3470 2740 3476
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2594 3431 2650 3440
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2792 2854 2820 3062
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2226 2000 2282 2009
rect 2226 1935 2282 1944
rect 2700 1601 2728 2790
rect 2884 2514 2912 3878
rect 2976 3194 3004 5034
rect 3068 4622 3096 5222
rect 3344 5080 3372 5578
rect 3436 5545 3464 5646
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3424 5092 3476 5098
rect 3344 5052 3424 5080
rect 3424 5034 3476 5040
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4859 3482 4868
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 4282 3096 4558
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3068 4049 3096 4082
rect 3054 4040 3110 4049
rect 3160 4010 3188 4490
rect 3436 4214 3464 4694
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3054 3975 3110 3984
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2976 2378 3004 2858
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2686 1592 2742 1601
rect 2686 1527 2742 1536
rect 2884 800 2912 2246
rect 3068 1970 3096 3538
rect 3344 3058 3372 3538
rect 3528 3534 3556 8230
rect 3606 7984 3662 7993
rect 3606 7919 3662 7928
rect 3620 7478 3648 7919
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3712 7342 3740 9046
rect 3790 8800 3846 8809
rect 3790 8735 3846 8744
rect 3804 7954 3832 8735
rect 3896 8537 3924 9646
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6458 3648 6598
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 6089 3648 6190
rect 3606 6080 3662 6089
rect 3606 6015 3662 6024
rect 3712 5658 3740 6802
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3620 5630 3740 5658
rect 3620 5370 3648 5630
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3712 5114 3740 5510
rect 3620 5086 3740 5114
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3422 3088 3478 3097
rect 3332 3052 3384 3058
rect 3422 3023 3424 3032
rect 3332 2994 3384 3000
rect 3476 3023 3478 3032
rect 3424 2994 3476 3000
rect 3620 2938 3648 5086
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3712 3058 3740 4966
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3620 2910 3740 2938
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 3620 2446 3648 2790
rect 3712 2582 3740 2910
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3056 1964 3108 1970
rect 3056 1906 3108 1912
rect 3712 800 3740 2246
rect 1674 776 1730 785
rect 1674 711 1730 720
rect 2042 0 2098 800
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 3804 377 3832 6598
rect 3896 5370 3924 8298
rect 3988 6934 4016 9522
rect 4080 9518 4108 11494
rect 4172 11393 4200 11562
rect 4158 11384 4214 11393
rect 4158 11319 4214 11328
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4172 9450 4200 11222
rect 4264 11218 4292 11562
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10266 4292 10950
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4356 10130 4384 10406
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4250 10024 4306 10033
rect 4250 9959 4252 9968
rect 4304 9959 4306 9968
rect 4252 9930 4304 9936
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4252 9580 4304 9586
rect 4356 9568 4384 9862
rect 4448 9654 4476 11648
rect 4528 11630 4580 11636
rect 4540 10810 4568 11630
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4540 10130 4568 10474
rect 4632 10441 4660 13382
rect 4894 13359 4950 13368
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 11694 4752 13262
rect 4908 12850 4936 13359
rect 5736 13326 5764 13631
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 5814 13424 5870 13433
rect 5814 13359 5870 13368
rect 6092 13388 6144 13394
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5828 13258 5856 13359
rect 6092 13330 6144 13336
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4908 12306 4936 12786
rect 5000 12753 5028 13126
rect 5092 12986 5120 13126
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 6012 12889 6040 13194
rect 5998 12880 6054 12889
rect 5632 12844 5684 12850
rect 5998 12815 6054 12824
rect 5632 12786 5684 12792
rect 4986 12744 5042 12753
rect 4986 12679 5042 12688
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4816 11354 4844 12038
rect 5000 11830 5028 12582
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5092 12238 5120 12378
rect 5644 12238 5672 12786
rect 6104 12714 6132 13330
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5092 11898 5120 12174
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5276 11898 5304 12038
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 5736 11898 5764 12038
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5828 11830 5856 12038
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 4986 11656 5042 11665
rect 4986 11591 5042 11600
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4908 10452 4936 11222
rect 5000 11121 5028 11591
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4986 11112 5042 11121
rect 4986 11047 5042 11056
rect 4988 11008 5040 11014
rect 4986 10976 4988 10985
rect 5040 10976 5042 10985
rect 4986 10911 5042 10920
rect 4986 10840 5042 10849
rect 4986 10775 4988 10784
rect 5040 10775 5042 10784
rect 4988 10746 5040 10752
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5000 10577 5028 10610
rect 5092 10606 5120 11494
rect 5828 11393 5856 11766
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5814 11384 5870 11393
rect 5814 11319 5870 11328
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5080 10600 5132 10606
rect 4986 10568 5042 10577
rect 5080 10542 5132 10548
rect 4986 10503 5042 10512
rect 4618 10432 4674 10441
rect 4908 10424 5120 10452
rect 5184 10441 5212 10610
rect 4618 10367 4674 10376
rect 4986 10296 5042 10305
rect 4986 10231 5042 10240
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4304 9540 4384 9568
rect 4252 9522 4304 9528
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4158 9344 4214 9353
rect 4158 9279 4214 9288
rect 4068 8832 4120 8838
rect 4172 8820 4200 9279
rect 4120 8792 4200 8820
rect 4068 8774 4120 8780
rect 4172 8673 4200 8792
rect 4158 8664 4214 8673
rect 4158 8599 4214 8608
rect 4172 8566 4200 8599
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4264 8242 4292 9522
rect 4540 9518 4568 10066
rect 4528 9512 4580 9518
rect 4526 9480 4528 9489
rect 4580 9480 4582 9489
rect 4344 9444 4396 9450
rect 4526 9415 4582 9424
rect 4344 9386 4396 9392
rect 4356 9024 4384 9386
rect 4632 9110 4660 10134
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4894 9888 4950 9897
rect 4816 9722 4844 9862
rect 4894 9823 4950 9832
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4804 9512 4856 9518
rect 4908 9500 4936 9823
rect 5000 9654 5028 10231
rect 5092 10062 5120 10424
rect 5170 10432 5226 10441
rect 5276 10418 5304 10950
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10843 5706 10852
rect 5814 10840 5870 10849
rect 5814 10775 5816 10784
rect 5868 10775 5870 10784
rect 5816 10746 5868 10752
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5448 10464 5500 10470
rect 5276 10390 5396 10418
rect 5448 10406 5500 10412
rect 5170 10367 5226 10376
rect 5262 10296 5318 10305
rect 5262 10231 5318 10240
rect 5276 10130 5304 10231
rect 5368 10198 5396 10390
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5080 10056 5132 10062
rect 5460 10033 5488 10406
rect 5644 10130 5672 10542
rect 5828 10146 5856 10610
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5736 10118 5856 10146
rect 5736 10033 5764 10118
rect 5080 9998 5132 10004
rect 5446 10024 5502 10033
rect 5446 9959 5502 9968
rect 5722 10024 5778 10033
rect 5722 9959 5778 9968
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5828 9586 5856 9930
rect 5920 9654 5948 11494
rect 6012 11218 6040 12582
rect 6288 11898 6316 13466
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12889 6408 13126
rect 6472 12918 6500 13670
rect 6826 13560 6882 13569
rect 6826 13495 6828 13504
rect 6880 13495 6882 13504
rect 6828 13466 6880 13472
rect 6840 13326 6868 13466
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6460 12912 6512 12918
rect 6366 12880 6422 12889
rect 6460 12854 6512 12860
rect 6366 12815 6422 12824
rect 6380 12782 6408 12815
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6564 12209 6592 13262
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6840 12730 6868 12922
rect 6748 12702 6868 12730
rect 6748 12646 6776 12702
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12238 6868 12582
rect 6828 12232 6880 12238
rect 6550 12200 6606 12209
rect 6828 12174 6880 12180
rect 6550 12135 6606 12144
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 9722 6040 10406
rect 6104 10062 6132 11630
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 4908 9472 5028 9500
rect 4804 9454 4856 9460
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4436 9036 4488 9042
rect 4356 8996 4436 9024
rect 4436 8978 4488 8984
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4448 8922 4476 8978
rect 4448 8894 4660 8922
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8634 4476 8774
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4080 8214 4292 8242
rect 4080 7449 4108 8214
rect 4356 8090 4384 8434
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4344 8084 4396 8090
rect 4172 8022 4200 8053
rect 4344 8026 4396 8032
rect 4160 8016 4212 8022
rect 4158 7984 4160 7993
rect 4212 7984 4214 7993
rect 4158 7919 4214 7928
rect 4252 7948 4304 7954
rect 4066 7440 4122 7449
rect 4172 7410 4200 7919
rect 4252 7890 4304 7896
rect 4066 7375 4122 7384
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3896 4826 3924 5102
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 2990 3924 4422
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3988 2922 4016 6734
rect 4080 4758 4108 7210
rect 4158 6760 4214 6769
rect 4158 6695 4160 6704
rect 4212 6695 4214 6704
rect 4160 6666 4212 6672
rect 4264 6440 4292 7890
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4342 7576 4398 7585
rect 4342 7511 4398 7520
rect 4356 7410 4384 7511
rect 4448 7449 4476 7754
rect 4434 7440 4490 7449
rect 4344 7404 4396 7410
rect 4434 7375 4490 7384
rect 4344 7346 4396 7352
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4172 6412 4292 6440
rect 4172 5681 4200 6412
rect 4356 6361 4384 6666
rect 4448 6390 4476 6734
rect 4436 6384 4488 6390
rect 4342 6352 4398 6361
rect 4252 6316 4304 6322
rect 4436 6326 4488 6332
rect 4342 6287 4398 6296
rect 4252 6258 4304 6264
rect 4264 5914 4292 6258
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4356 5953 4384 6190
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4342 5944 4398 5953
rect 4252 5908 4304 5914
rect 4342 5879 4398 5888
rect 4252 5850 4304 5856
rect 4158 5672 4214 5681
rect 4158 5607 4214 5616
rect 4172 5098 4200 5607
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3882 2680 3938 2689
rect 3882 2615 3884 2624
rect 3936 2615 3938 2624
rect 3884 2586 3936 2592
rect 4080 2514 4108 4422
rect 4172 3738 4200 4558
rect 4264 4026 4292 5850
rect 4448 5658 4476 6054
rect 4540 5778 4568 8366
rect 4632 7698 4660 8894
rect 4724 7954 4752 8978
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4816 7886 4844 9454
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8906 4936 9318
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4632 7670 4936 7698
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4632 5778 4660 7142
rect 4724 6202 4752 7278
rect 4724 6174 4844 6202
rect 4712 6112 4764 6118
rect 4816 6089 4844 6174
rect 4712 6054 4764 6060
rect 4802 6080 4858 6089
rect 4724 5817 4752 6054
rect 4802 6015 4858 6024
rect 4804 5840 4856 5846
rect 4710 5808 4766 5817
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4620 5772 4672 5778
rect 4804 5782 4856 5788
rect 4710 5743 4766 5752
rect 4620 5714 4672 5720
rect 4712 5704 4764 5710
rect 4448 5630 4660 5658
rect 4712 5646 4764 5652
rect 4632 5574 4660 5630
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4448 4264 4476 5510
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4356 4236 4476 4264
rect 4356 4128 4384 4236
rect 4540 4214 4568 4762
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4356 4100 4476 4128
rect 4264 3998 4384 4026
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 3194 4292 3878
rect 4356 3534 4384 3998
rect 4448 3602 4476 4100
rect 4540 3602 4568 4150
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4344 3392 4396 3398
rect 4342 3360 4344 3369
rect 4528 3392 4580 3398
rect 4396 3360 4398 3369
rect 4528 3334 4580 3340
rect 4342 3295 4398 3304
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4356 2961 4384 3295
rect 4342 2952 4398 2961
rect 4342 2887 4398 2896
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4540 800 4568 3334
rect 4632 3194 4660 5034
rect 4724 4486 4752 5646
rect 4816 5370 4844 5782
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4908 5250 4936 7670
rect 5000 6304 5028 9472
rect 5920 9450 6040 9466
rect 5920 9444 6052 9450
rect 5920 9438 6000 9444
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 7857 5120 8774
rect 5184 7954 5212 9318
rect 5920 9217 5948 9438
rect 6000 9386 6052 9392
rect 5998 9344 6054 9353
rect 5998 9279 6054 9288
rect 5906 9208 5962 9217
rect 5906 9143 5962 9152
rect 5630 9072 5686 9081
rect 5630 9007 5632 9016
rect 5684 9007 5686 9016
rect 5632 8978 5684 8984
rect 5816 8968 5868 8974
rect 5814 8936 5816 8945
rect 5868 8936 5870 8945
rect 5814 8871 5870 8880
rect 5920 8838 5948 9143
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 5736 8090 5764 8774
rect 5920 8430 5948 8774
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5264 7880 5316 7886
rect 5078 7848 5134 7857
rect 5724 7880 5776 7886
rect 5264 7822 5316 7828
rect 5722 7848 5724 7857
rect 5776 7848 5778 7857
rect 5078 7783 5134 7792
rect 5276 7546 5304 7822
rect 5828 7818 5856 8298
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 8090 5948 8230
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5722 7783 5778 7792
rect 5816 7812 5868 7818
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5080 6316 5132 6322
rect 5000 6276 5080 6304
rect 5080 6258 5132 6264
rect 5184 6118 5212 7278
rect 5276 6730 5304 7482
rect 5538 7440 5594 7449
rect 5538 7375 5540 7384
rect 5592 7375 5594 7384
rect 5540 7346 5592 7352
rect 5736 6905 5764 7783
rect 5816 7754 5868 7760
rect 5920 7274 5948 7822
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5722 6896 5778 6905
rect 5722 6831 5778 6840
rect 5920 6798 5948 7210
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5724 6656 5776 6662
rect 5776 6604 5856 6610
rect 5724 6598 5856 6604
rect 5736 6582 5856 6598
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 5828 6322 5856 6582
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5953 5212 6054
rect 5170 5944 5226 5953
rect 5170 5879 5226 5888
rect 5368 5846 5396 6258
rect 5814 6216 5870 6225
rect 5814 6151 5870 6160
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5828 5778 5856 6151
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4816 5222 4936 5250
rect 4816 4826 4844 5222
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4712 4140 4764 4146
rect 4764 4100 4844 4128
rect 4712 4082 4764 4088
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4724 3738 4752 3946
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4724 2938 4752 3402
rect 4816 3058 4844 4100
rect 4908 3466 4936 5102
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4632 2378 4660 2926
rect 4724 2910 4936 2938
rect 5000 2922 5028 5510
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5080 5160 5132 5166
rect 5132 5108 5212 5114
rect 5080 5102 5212 5108
rect 5092 5086 5212 5102
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5092 4146 5120 4558
rect 5184 4486 5212 5086
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5092 3194 5120 4082
rect 5184 3398 5212 4422
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5276 3074 5304 5170
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5460 4622 5488 5034
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 5736 4282 5764 5102
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5908 4140 5960 4146
rect 5828 4100 5908 4128
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3534 5764 3878
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 5828 3126 5856 4100
rect 5908 4082 5960 4088
rect 5184 3046 5304 3074
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5184 2990 5212 3046
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4802 2816 4858 2825
rect 4724 2582 4752 2790
rect 4802 2751 4858 2760
rect 4908 2774 4936 2910
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4816 2446 4844 2751
rect 4908 2746 5028 2774
rect 5000 2514 5028 2746
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4632 2106 4660 2314
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 5276 1170 5304 2586
rect 6012 2446 6040 9279
rect 6104 8498 6132 9998
rect 6196 9926 6224 10610
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6288 9518 6316 11154
rect 6380 10810 6408 11494
rect 6564 11234 6592 11562
rect 6656 11354 6684 11698
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6564 11206 6684 11234
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6380 10441 6408 10746
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6366 10432 6422 10441
rect 6366 10367 6422 10376
rect 6380 10266 6408 10367
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9722 6408 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6104 4826 6132 8434
rect 6196 8294 6224 9454
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6380 9353 6408 9386
rect 6472 9382 6500 10542
rect 6460 9376 6512 9382
rect 6366 9344 6422 9353
rect 6460 9318 6512 9324
rect 6366 9279 6422 9288
rect 6564 9194 6592 11018
rect 6656 10996 6684 11206
rect 6748 11150 6776 11630
rect 6932 11626 6960 13330
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12918 7052 13126
rect 7392 12986 7420 13903
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7392 12434 7420 12718
rect 7300 12406 7420 12434
rect 7300 12238 7328 12406
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11150 6868 11494
rect 7024 11218 7052 12038
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7116 11762 7144 11834
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6736 11144 6788 11150
rect 6828 11144 6880 11150
rect 6736 11086 6788 11092
rect 6826 11112 6828 11121
rect 6880 11112 6882 11121
rect 6826 11047 6882 11056
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6656 10968 6776 10996
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9761 6684 10066
rect 6642 9752 6698 9761
rect 6642 9687 6698 9696
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6380 9166 6592 9194
rect 6274 9072 6330 9081
rect 6274 9007 6330 9016
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6288 6662 6316 9007
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6196 6118 6224 6258
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6288 5302 6316 6598
rect 6380 6322 6408 9166
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6288 4729 6316 4966
rect 6274 4720 6330 4729
rect 6274 4655 6330 4664
rect 6380 4554 6408 6054
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6196 3126 6224 3470
rect 6184 3120 6236 3126
rect 6090 3088 6146 3097
rect 6184 3062 6236 3068
rect 6090 3023 6092 3032
rect 6144 3023 6146 3032
rect 6092 2994 6144 3000
rect 6196 2990 6224 3062
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6288 2774 6316 3878
rect 6196 2746 6316 2774
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 5276 1142 5396 1170
rect 5368 800 5396 1142
rect 6196 800 6224 2746
rect 6472 2446 6500 9046
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8566 6592 8910
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6656 8430 6684 9522
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6550 8256 6606 8265
rect 6550 8191 6606 8200
rect 6564 6118 6592 8191
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6656 6254 6684 7346
rect 6748 7324 6776 10968
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 9897 6868 10542
rect 6826 9888 6882 9897
rect 6826 9823 6882 9832
rect 6932 9738 6960 11018
rect 7024 10606 7052 11154
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10198 7052 10406
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6932 9710 7052 9738
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 8906 6868 9454
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6840 8634 6868 8842
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6932 7478 6960 9318
rect 7024 7818 7052 9710
rect 7116 9500 7144 11562
rect 7208 11121 7236 12038
rect 7194 11112 7250 11121
rect 7300 11082 7328 12174
rect 7194 11047 7250 11056
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 9926 7236 10950
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7196 9512 7248 9518
rect 7116 9472 7196 9500
rect 7196 9454 7248 9460
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8022 7144 8774
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6748 7296 6960 7324
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6254 6868 7142
rect 6932 6882 6960 7296
rect 7024 7002 7052 7754
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6932 6854 7052 6882
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5704 6696 5710
rect 6748 5681 6776 6054
rect 6840 5710 6868 6190
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5704 6880 5710
rect 6644 5646 6696 5652
rect 6734 5672 6790 5681
rect 6656 5234 6684 5646
rect 6828 5646 6880 5652
rect 6734 5607 6790 5616
rect 6748 5273 6776 5607
rect 6734 5264 6790 5273
rect 6644 5228 6696 5234
rect 6734 5199 6790 5208
rect 6644 5170 6696 5176
rect 6656 4808 6684 5170
rect 6828 4820 6880 4826
rect 6656 4780 6828 4808
rect 6656 4622 6684 4780
rect 6828 4762 6880 4768
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6932 4185 6960 6054
rect 7024 5522 7052 6854
rect 7116 5642 7144 7958
rect 7208 6662 7236 9454
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7024 5494 7236 5522
rect 7208 5234 7236 5494
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7102 5128 7158 5137
rect 7102 5063 7158 5072
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 6918 4176 6974 4185
rect 6552 4140 6604 4146
rect 6918 4111 6974 4120
rect 6552 4082 6604 4088
rect 6564 3670 6592 4082
rect 7024 4010 7052 4490
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 7116 3058 7144 5063
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7208 2854 7236 5170
rect 7300 4554 7328 10066
rect 7392 8480 7420 12242
rect 7484 11286 7512 12718
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 8128 12434 8156 14282
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 7944 12406 8156 12434
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11898 7696 12038
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 11626 7788 11834
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7944 11558 7972 12406
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7576 11150 7604 11290
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7668 10606 7696 11154
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 10062 7512 10406
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 8036 10266 8064 10474
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7470 9888 7526 9897
rect 7470 9823 7526 9832
rect 7484 9092 7512 9823
rect 7852 9625 7880 10134
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7944 9761 7972 9862
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 7838 9616 7894 9625
rect 7838 9551 7894 9560
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 8036 9178 8064 9522
rect 8128 9450 8156 12174
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11898 8524 12038
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11150 8432 11494
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8588 11218 8616 11290
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8772 11082 8800 11630
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10198 8248 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8220 9450 8248 9930
rect 8312 9722 8340 9930
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8312 9178 8340 9454
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 7484 9064 7604 9092
rect 7472 8492 7524 8498
rect 7392 8452 7472 8480
rect 7392 8090 7420 8452
rect 7472 8434 7524 8440
rect 7576 8378 7604 9064
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8022 8392 8078 8401
rect 7484 8350 7604 8378
rect 7944 8350 8022 8378
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7392 7410 7420 7686
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7378 6080 7434 6089
rect 7378 6015 7434 6024
rect 7392 5302 7420 6015
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 7300 2378 7328 4490
rect 7484 4486 7512 8350
rect 7944 8294 7972 8350
rect 8022 8327 8078 8336
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 7206 7604 7890
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4859 7930 4868
rect 8036 4826 8064 8327
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5234 8156 5646
rect 8220 5574 8248 8774
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 6118 8340 6666
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 8036 3482 8064 4150
rect 8404 4146 8432 10066
rect 8496 7546 8524 11018
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8588 9654 8616 10542
rect 8680 10062 8708 10542
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8666 9616 8722 9625
rect 8666 9551 8722 9560
rect 8576 9512 8628 9518
rect 8680 9500 8708 9551
rect 8628 9472 8708 9500
rect 8576 9454 8628 9460
rect 8588 9081 8616 9454
rect 8574 9072 8630 9081
rect 8574 9007 8630 9016
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 7944 3454 8064 3482
rect 8128 3466 8156 3946
rect 8220 3602 8248 4082
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8116 3460 8168 3466
rect 7944 3398 7972 3454
rect 8116 3402 8168 3408
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6564 2038 6592 2246
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6932 1170 6960 2246
rect 7392 2106 7420 2314
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7944 1970 7972 2246
rect 7932 1964 7984 1970
rect 7932 1906 7984 1912
rect 6932 1142 7052 1170
rect 7024 800 7052 1142
rect 8036 898 8064 3334
rect 8220 3126 8248 3538
rect 8496 3534 8524 7482
rect 8680 6798 8708 8978
rect 8772 7750 8800 11018
rect 8956 11014 8984 13806
rect 9586 13288 9642 13297
rect 9586 13223 9642 13232
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12102 9260 12650
rect 9324 12238 9352 12718
rect 9600 12434 9628 13223
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12442 9720 12582
rect 9508 12406 9628 12434
rect 9680 12436 9732 12442
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9402 12064 9458 12073
rect 9232 11830 9260 12038
rect 9402 11999 9458 12008
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9220 11688 9272 11694
rect 9218 11656 9220 11665
rect 9272 11656 9274 11665
rect 9218 11591 9274 11600
rect 9232 11121 9260 11591
rect 9324 11558 9352 11698
rect 9416 11665 9444 11999
rect 9508 11830 9536 12406
rect 10244 12434 10272 14214
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13841 10548 13874
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10888 13734 10916 14350
rect 12820 14074 12848 14350
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13832 13938 13860 14350
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 9732 12406 9812 12434
rect 10244 12406 10364 12434
rect 9680 12378 9732 12384
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9692 11830 9720 12271
rect 9784 12238 9812 12406
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10244 12238 10272 12310
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 11898 9812 12038
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9496 11688 9548 11694
rect 9402 11656 9458 11665
rect 9496 11630 9548 11636
rect 9402 11591 9458 11600
rect 9312 11552 9364 11558
rect 9310 11520 9312 11529
rect 9364 11520 9366 11529
rect 9310 11455 9366 11464
rect 9324 11429 9352 11455
rect 9218 11112 9274 11121
rect 9218 11047 9274 11056
rect 9232 11014 9260 11047
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8864 9926 8892 10746
rect 8956 10470 8984 10950
rect 9034 10840 9090 10849
rect 9034 10775 9090 10784
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8956 9722 8984 10066
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9048 9674 9076 10775
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9324 9722 9352 10134
rect 9312 9716 9364 9722
rect 9048 9646 9260 9674
rect 9312 9658 9364 9664
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8864 7886 8892 8502
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8864 7478 8892 7822
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8864 6866 8892 7414
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8956 6662 8984 9454
rect 9048 8362 9076 9646
rect 9232 9586 9260 9646
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9140 8786 9168 9522
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9232 8906 9260 9386
rect 9324 9110 9352 9658
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9140 8758 9260 8786
rect 9232 8498 9260 8758
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 8022 9076 8298
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9232 6730 9260 8434
rect 9324 7993 9352 8842
rect 9416 8838 9444 9114
rect 9508 9042 9536 11630
rect 9600 11150 9628 11698
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9680 11144 9732 11150
rect 9876 11132 9904 11494
rect 9732 11104 9904 11132
rect 10152 11132 10180 11630
rect 10244 11257 10272 12174
rect 10230 11248 10286 11257
rect 10230 11183 10286 11192
rect 10152 11104 10272 11132
rect 9680 11086 9732 11092
rect 9600 10130 9628 11086
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 10244 10810 10272 11104
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8294 9444 8774
rect 9494 8528 9550 8537
rect 9494 8463 9550 8472
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9404 7404 9456 7410
rect 9508 7392 9536 8463
rect 9456 7364 9536 7392
rect 9404 7346 9456 7352
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6322 8984 6598
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5710 9260 6190
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9324 5370 9352 5578
rect 9416 5370 9444 7346
rect 9496 6316 9548 6322
rect 9548 6276 9628 6304
rect 9496 6258 9548 6264
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9600 5030 9628 6276
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 8772 3942 8800 4966
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8404 3058 8432 3334
rect 8588 3058 8616 3674
rect 9402 3632 9458 3641
rect 9402 3567 9458 3576
rect 9416 3534 9444 3567
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8116 2984 8168 2990
rect 8114 2952 8116 2961
rect 8300 2984 8352 2990
rect 8168 2952 8170 2961
rect 8300 2926 8352 2932
rect 8114 2887 8170 2896
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8128 1970 8156 2790
rect 8312 2446 8340 2926
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8116 1964 8168 1970
rect 8116 1906 8168 1912
rect 7852 870 8064 898
rect 7852 800 7880 870
rect 8680 800 8708 2790
rect 8772 2446 8800 3334
rect 9140 2650 9168 3470
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9324 3194 9352 3402
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9232 2378 9260 2790
rect 9600 2650 9628 4490
rect 9692 2854 9720 9454
rect 9784 9178 9812 10610
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 9846 9820 10154 9829
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 10244 9722 10272 10406
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10230 9480 10286 9489
rect 9968 9178 9996 9454
rect 10230 9415 10286 9424
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9864 9036 9916 9042
rect 9784 8974 9812 9007
rect 10048 9036 10100 9042
rect 9916 8996 10048 9024
rect 9864 8978 9916 8984
rect 10048 8978 10100 8984
rect 10152 8974 10180 9318
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9864 8832 9916 8838
rect 9784 8792 9864 8820
rect 9784 3534 9812 8792
rect 9864 8774 9916 8780
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 10244 8634 10272 9415
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10244 7993 10272 8570
rect 10230 7984 10286 7993
rect 10230 7919 10286 7928
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 10244 7002 10272 7754
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10244 5710 10272 6190
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5403 10154 5412
rect 10336 5250 10364 12406
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10428 12170 10456 12310
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10414 12064 10470 12073
rect 10414 11999 10470 12008
rect 10428 11626 10456 11999
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10416 11280 10468 11286
rect 10414 11248 10416 11257
rect 10468 11248 10470 11257
rect 10414 11183 10470 11192
rect 10520 11150 10548 11494
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10612 11098 10640 12786
rect 10782 11656 10838 11665
rect 10782 11591 10838 11600
rect 10612 11070 10732 11098
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10428 9450 10456 10542
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10520 9382 10548 9862
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10244 5234 10364 5250
rect 10232 5228 10364 5234
rect 10284 5222 10364 5228
rect 10232 5170 10284 5176
rect 10138 4720 10194 4729
rect 10138 4655 10194 4664
rect 10152 4622 10180 4655
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 10428 3754 10456 7822
rect 10612 7818 10640 10950
rect 10704 10130 10732 11070
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10796 9704 10824 11591
rect 10704 9676 10824 9704
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10704 7274 10732 9676
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10704 6322 10732 7210
rect 10796 6662 10824 9454
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10598 5672 10654 5681
rect 10704 5642 10732 6054
rect 10598 5607 10654 5616
rect 10692 5636 10744 5642
rect 10612 4622 10640 5607
rect 10692 5578 10744 5584
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10612 4185 10640 4558
rect 10598 4176 10654 4185
rect 10598 4111 10654 4120
rect 10336 3726 10456 3754
rect 10336 3670 10364 3726
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9772 3392 9824 3398
rect 10336 3380 10364 3606
rect 9772 3334 9824 3340
rect 10244 3352 10364 3380
rect 9784 3194 9812 3334
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 10244 3058 10272 3352
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9496 2576 9548 2582
rect 9402 2544 9458 2553
rect 9496 2518 9548 2524
rect 9402 2479 9458 2488
rect 9416 2378 9444 2479
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9508 800 9536 2518
rect 10060 2446 10088 2994
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 1902 9812 2246
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 10336 800 10364 2790
rect 10704 2310 10732 5170
rect 10888 3398 10916 13670
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12434 11192 13126
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 11794 12744 11850 12753
rect 11794 12679 11850 12688
rect 11164 12406 11468 12434
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 11694 11008 12242
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11014 11008 11630
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10980 10470 11008 10610
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10266 11008 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 4593 11008 10066
rect 10966 4584 11022 4593
rect 10966 4519 11022 4528
rect 11072 3738 11100 11290
rect 11256 11218 11284 11562
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11256 10690 11284 11154
rect 11164 10662 11284 10690
rect 11334 10704 11390 10713
rect 11164 8566 11192 10662
rect 11334 10639 11336 10648
rect 11388 10639 11390 10648
rect 11336 10610 11388 10616
rect 11440 10169 11468 12406
rect 11808 12102 11836 12679
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 12530 12472 12586 12481
rect 12530 12407 12532 12416
rect 12584 12407 12586 12416
rect 12532 12378 12584 12384
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11808 11801 11836 12038
rect 11992 11898 12020 12038
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11794 11792 11850 11801
rect 11794 11727 11850 11736
rect 12084 11694 12112 12242
rect 12452 11830 12480 12310
rect 12636 12102 12664 12786
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11532 10198 11560 11018
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11702 10704 11758 10713
rect 11702 10639 11758 10648
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11520 10192 11572 10198
rect 11426 10160 11482 10169
rect 11520 10134 11572 10140
rect 11426 10095 11482 10104
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9722 11284 9862
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11348 9081 11376 9998
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11334 9072 11390 9081
rect 11244 9036 11296 9042
rect 11334 9007 11336 9016
rect 11244 8978 11296 8984
rect 11388 9007 11390 9016
rect 11336 8978 11388 8984
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11164 6730 11192 8502
rect 11256 7886 11284 8978
rect 11348 8947 11376 8978
rect 11440 8838 11468 9318
rect 11532 9178 11560 10134
rect 11624 9382 11652 10542
rect 11716 10033 11744 10639
rect 11808 10470 11836 10950
rect 11992 10742 12020 11630
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 11980 10736 12032 10742
rect 11900 10696 11980 10724
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11702 10024 11758 10033
rect 11702 9959 11758 9968
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11520 9036 11572 9042
rect 11624 9024 11652 9318
rect 11808 9081 11836 10406
rect 11900 10198 11928 10696
rect 11980 10678 12032 10684
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11888 10056 11940 10062
rect 11886 10024 11888 10033
rect 11940 10024 11942 10033
rect 11886 9959 11942 9968
rect 11572 8996 11652 9024
rect 11794 9072 11850 9081
rect 11794 9007 11850 9016
rect 11520 8978 11572 8984
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11348 7954 11376 8434
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7206 11284 7686
rect 11348 7410 11376 7890
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5273 11192 6054
rect 11150 5264 11206 5273
rect 11150 5199 11206 5208
rect 11164 4049 11192 5199
rect 11256 4146 11284 7142
rect 11348 6866 11376 7346
rect 11440 7002 11468 7822
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11348 5710 11376 6802
rect 11532 6254 11560 8978
rect 11610 8392 11666 8401
rect 11610 8327 11666 8336
rect 11624 7410 11652 8327
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11702 7304 11758 7313
rect 11702 7239 11758 7248
rect 11716 6633 11744 7239
rect 11702 6624 11758 6633
rect 11702 6559 11758 6568
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11624 5778 11652 6122
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11348 5302 11376 5646
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11348 4690 11376 5238
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4826 11468 4966
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11348 4214 11376 4626
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11150 4040 11206 4049
rect 11150 3975 11206 3984
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11256 3505 11284 3878
rect 11348 3602 11376 4150
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11242 3496 11298 3505
rect 11242 3431 11298 3440
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 11348 3126 11376 3538
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 11164 800 11192 2858
rect 11348 2514 11376 3062
rect 11440 2854 11468 4082
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11532 2650 11560 4490
rect 11624 4010 11652 5714
rect 11716 5681 11744 6054
rect 11702 5672 11758 5681
rect 11702 5607 11758 5616
rect 11808 5522 11836 9007
rect 11716 5494 11836 5522
rect 11716 4146 11744 5494
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11808 4282 11836 4558
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11900 4146 11928 9959
rect 11992 9722 12020 10406
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 12452 10169 12480 10542
rect 12636 10470 12664 10746
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 10192 12584 10198
rect 12438 10160 12494 10169
rect 12072 10124 12124 10130
rect 12532 10134 12584 10140
rect 12438 10095 12494 10104
rect 12072 10066 12124 10072
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 12084 9518 12112 10066
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12072 9512 12124 9518
rect 11992 9472 12072 9500
rect 11992 6730 12020 9472
rect 12072 9454 12124 9460
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 12452 9042 12480 9522
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 12452 6769 12480 8570
rect 12162 6760 12218 6769
rect 11980 6724 12032 6730
rect 12162 6695 12218 6704
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 11980 6666 12032 6672
rect 11992 5794 12020 6666
rect 12176 6361 12204 6695
rect 12438 6624 12494 6633
rect 12438 6559 12494 6568
rect 12254 6488 12310 6497
rect 12452 6458 12480 6559
rect 12254 6423 12256 6432
rect 12308 6423 12310 6432
rect 12440 6452 12492 6458
rect 12256 6394 12308 6400
rect 12440 6394 12492 6400
rect 12162 6352 12218 6361
rect 12162 6287 12218 6296
rect 12176 6254 12204 6287
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12072 5840 12124 5846
rect 11992 5788 12072 5794
rect 11992 5782 12124 5788
rect 12254 5808 12310 5817
rect 11992 5766 12112 5782
rect 12254 5743 12256 5752
rect 12308 5743 12310 5752
rect 12256 5714 12308 5720
rect 12360 5574 12388 5850
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11992 5030 12020 5306
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11992 3534 12020 4966
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4859 12378 4868
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12268 4282 12296 4490
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 12360 3942 12388 3975
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12360 3466 12388 3606
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 3194 11836 3334
rect 12452 3194 12480 4422
rect 12544 3602 12572 10134
rect 12636 9994 12664 10406
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12728 9874 12756 11630
rect 12912 10810 12940 13874
rect 13544 13864 13596 13870
rect 13542 13832 13544 13841
rect 14004 13864 14056 13870
rect 13596 13832 13598 13841
rect 14004 13806 14056 13812
rect 13542 13767 13598 13776
rect 13450 13288 13506 13297
rect 13268 13252 13320 13258
rect 13450 13223 13506 13232
rect 13268 13194 13320 13200
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12238 13032 12582
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11150 13124 11494
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13188 10690 13216 11086
rect 12912 10662 13216 10690
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 10130 12848 10474
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12636 9846 12756 9874
rect 12636 9518 12664 9846
rect 12820 9654 12848 10066
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12636 8838 12664 9046
rect 12820 9042 12848 9454
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 6118 12664 8774
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12636 2961 12664 6054
rect 12728 4146 12756 8298
rect 12820 6882 12848 8978
rect 12912 7834 12940 10662
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13004 8362 13032 10066
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9722 13124 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12990 7848 13046 7857
rect 12912 7806 12990 7834
rect 12990 7783 13046 7792
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12912 7449 12940 7482
rect 12898 7440 12954 7449
rect 12898 7375 12954 7384
rect 13004 7342 13032 7783
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12990 6896 13046 6905
rect 12820 6854 12990 6882
rect 12990 6831 12992 6840
rect 13044 6831 13046 6840
rect 12992 6802 13044 6808
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12806 6352 12862 6361
rect 12912 6322 12940 6598
rect 13004 6497 13032 6802
rect 12990 6488 13046 6497
rect 12990 6423 13046 6432
rect 12806 6287 12808 6296
rect 12860 6287 12862 6296
rect 12900 6316 12952 6322
rect 12808 6258 12860 6264
rect 12900 6258 12952 6264
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12912 3534 12940 6054
rect 13004 3534 13032 6190
rect 13096 5642 13124 9454
rect 13188 8362 13216 10474
rect 13280 9568 13308 13194
rect 13464 12918 13492 13223
rect 13452 12912 13504 12918
rect 13450 12880 13452 12889
rect 13504 12880 13506 12889
rect 13450 12815 13506 12824
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12442 13768 12582
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13360 12096 13412 12102
rect 13464 12084 13492 12378
rect 14016 12322 14044 13806
rect 14108 13025 14136 14214
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 15212 13734 15240 14282
rect 15304 13802 15332 14894
rect 15476 14544 15528 14550
rect 15474 14512 15476 14521
rect 15528 14512 15530 14521
rect 15474 14447 15530 14456
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14094 13016 14150 13025
rect 14294 13019 14602 13028
rect 14094 12951 14150 12960
rect 14108 12374 14136 12951
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14554 12472 14610 12481
rect 14554 12407 14610 12416
rect 13648 12294 14044 12322
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 13412 12056 13492 12084
rect 13544 12096 13596 12102
rect 13360 12038 13412 12044
rect 13544 12038 13596 12044
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13464 11218 13492 11698
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13464 10810 13492 10950
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13372 9722 13400 9998
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13280 9540 13400 9568
rect 13266 9480 13322 9489
rect 13266 9415 13322 9424
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13188 6458 13216 8298
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13280 5914 13308 9415
rect 13372 9092 13400 9540
rect 13464 9217 13492 10542
rect 13556 10062 13584 12038
rect 13648 11762 13676 12294
rect 14568 12238 14596 12407
rect 14660 12306 14688 12718
rect 14844 12434 14872 13126
rect 15120 12481 15148 13262
rect 15396 13258 15424 14350
rect 15672 14006 15700 14418
rect 16040 14346 16068 16079
rect 16210 15736 16266 15745
rect 16210 15671 16266 15680
rect 16224 14822 16252 15671
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14346 16252 14758
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16040 14226 16068 14282
rect 15948 14198 16068 14226
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15948 13938 15976 14198
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16028 13932 16080 13938
rect 16132 13920 16160 14214
rect 16316 13938 16344 16487
rect 16578 16400 16634 16510
rect 16394 15328 16450 15337
rect 16394 15263 16450 15272
rect 16408 14414 16436 15263
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 16868 14482 16896 16510
rect 18786 16400 18842 17200
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16396 14408 16448 14414
rect 17040 14408 17092 14414
rect 16396 14350 16448 14356
rect 16670 14376 16726 14385
rect 17040 14350 17092 14356
rect 16670 14311 16726 14320
rect 16684 13938 16712 14311
rect 16080 13892 16160 13920
rect 16304 13932 16356 13938
rect 16028 13874 16080 13880
rect 16304 13874 16356 13880
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 15488 13841 15516 13874
rect 15474 13832 15530 13841
rect 16854 13832 16910 13841
rect 15474 13767 15530 13776
rect 16120 13796 16172 13802
rect 16854 13767 16856 13776
rect 16120 13738 16172 13744
rect 16908 13767 16910 13776
rect 16856 13738 16908 13744
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 14752 12406 14872 12434
rect 15106 12472 15162 12481
rect 15106 12407 15162 12416
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 13912 12232 13964 12238
rect 13818 12200 13874 12209
rect 13912 12174 13964 12180
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 13818 12135 13874 12144
rect 13832 12102 13860 12135
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 11937 13860 12038
rect 13818 11928 13874 11937
rect 13818 11863 13874 11872
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11218 13768 11630
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13648 9654 13676 10678
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13450 9208 13506 9217
rect 13450 9143 13506 9152
rect 13372 9064 13492 9092
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13372 8537 13400 8570
rect 13358 8528 13414 8537
rect 13358 8463 13414 8472
rect 13464 7206 13492 9064
rect 13556 9042 13584 9522
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9110 13676 9454
rect 13740 9382 13768 11018
rect 13832 10742 13860 11018
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8673 13676 8910
rect 13634 8664 13690 8673
rect 13740 8634 13768 9318
rect 13634 8599 13690 8608
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 7880 13688 7886
rect 13634 7848 13636 7857
rect 13688 7848 13690 7857
rect 13634 7783 13690 7792
rect 13648 7585 13676 7783
rect 13634 7576 13690 7585
rect 13832 7546 13860 10542
rect 13924 10130 13952 12174
rect 14016 12102 14044 12174
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14200 11830 14228 12106
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14568 11626 14596 11766
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11150 14412 11494
rect 14568 11257 14596 11562
rect 14554 11248 14610 11257
rect 14554 11183 14610 11192
rect 14372 11144 14424 11150
rect 14094 11112 14150 11121
rect 14372 11086 14424 11092
rect 14094 11047 14150 11056
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 14016 9761 14044 10406
rect 14002 9752 14058 9761
rect 13912 9716 13964 9722
rect 14002 9687 14058 9696
rect 13912 9658 13964 9664
rect 13634 7511 13690 7520
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13544 7336 13596 7342
rect 13542 7304 13544 7313
rect 13596 7304 13598 7313
rect 13542 7239 13598 7248
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13740 6798 13768 6870
rect 13728 6792 13780 6798
rect 13634 6760 13690 6769
rect 13728 6734 13780 6740
rect 13634 6695 13690 6704
rect 13648 6662 13676 6695
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13636 6656 13688 6662
rect 13740 6633 13768 6734
rect 13636 6598 13688 6604
rect 13726 6624 13782 6633
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4282 13124 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12622 2952 12678 2961
rect 12622 2887 12678 2896
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11992 800 12020 2586
rect 12728 1834 12756 3334
rect 12716 1828 12768 1834
rect 12716 1770 12768 1776
rect 12820 800 12848 3334
rect 13096 2446 13124 3402
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13188 2582 13216 2790
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 2514 13308 2994
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13004 2038 13032 2382
rect 13372 2038 13400 6598
rect 13726 6559 13782 6568
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 5234 13768 5510
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3602 13584 4082
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13464 3194 13492 3402
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13556 3058 13584 3538
rect 13740 3126 13768 4694
rect 13832 4078 13860 7482
rect 13924 5710 13952 9658
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14016 8129 14044 9590
rect 14002 8120 14058 8129
rect 14002 8055 14058 8064
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3126 13860 3878
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13820 3120 13872 3126
rect 14016 3097 14044 7686
rect 14108 7410 14136 11047
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 9382 14228 10610
rect 14660 10606 14688 12242
rect 14752 11558 14780 12406
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 15014 12336 15070 12345
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14738 10840 14794 10849
rect 14738 10775 14794 10784
rect 14752 10742 14780 10775
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10062 14504 10406
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 14738 9752 14794 9761
rect 14648 9716 14700 9722
rect 14700 9696 14738 9704
rect 14700 9687 14794 9696
rect 14700 9676 14780 9687
rect 14648 9658 14700 9664
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14370 9344 14426 9353
rect 14370 9279 14426 9288
rect 14186 9208 14242 9217
rect 14186 9143 14242 9152
rect 14200 7528 14228 9143
rect 14384 8838 14412 9279
rect 14462 9208 14518 9217
rect 14568 9178 14596 9386
rect 14844 9353 14872 12310
rect 15014 12271 15070 12280
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14936 11286 14964 11698
rect 15028 11354 15056 12271
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 14936 9654 14964 11222
rect 15028 11098 15056 11290
rect 15028 11070 15240 11098
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10810 15148 10950
rect 15212 10810 15240 11070
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15212 10554 15240 10746
rect 15212 10526 15332 10554
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15028 9722 15056 9862
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14924 9376 14976 9382
rect 14830 9344 14886 9353
rect 14924 9318 14976 9324
rect 14830 9279 14886 9288
rect 14936 9194 14964 9318
rect 14462 9143 14518 9152
rect 14556 9172 14608 9178
rect 14476 9110 14504 9143
rect 14556 9114 14608 9120
rect 14660 9166 14964 9194
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14556 9036 14608 9042
rect 14660 9024 14688 9166
rect 14924 9104 14976 9110
rect 14608 8996 14688 9024
rect 14830 9072 14886 9081
rect 14924 9046 14976 9052
rect 14830 9007 14832 9016
rect 14556 8978 14608 8984
rect 14884 9007 14886 9016
rect 14832 8978 14884 8984
rect 14936 8838 14964 9046
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 14752 8673 14780 8774
rect 14738 8664 14794 8673
rect 14738 8599 14794 8608
rect 15028 8514 15056 8978
rect 14844 8498 15056 8514
rect 14832 8492 15056 8498
rect 14884 8486 15056 8492
rect 14832 8434 14884 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14476 8022 14504 8366
rect 15120 8294 15148 10066
rect 15212 9586 15240 10406
rect 15304 9897 15332 10526
rect 15396 10062 15424 11290
rect 15488 11150 15516 11494
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15488 10130 15516 10542
rect 15580 10305 15608 11154
rect 15566 10296 15622 10305
rect 15566 10231 15622 10240
rect 15580 10130 15608 10231
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15384 9920 15436 9926
rect 15290 9888 15346 9897
rect 15384 9862 15436 9868
rect 15290 9823 15346 9832
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15212 9178 15240 9522
rect 15304 9178 15332 9590
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15212 9058 15240 9114
rect 15212 9030 15332 9058
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15212 8809 15240 8910
rect 15198 8800 15254 8809
rect 15198 8735 15254 8744
rect 15304 8566 15332 9030
rect 15396 8838 15424 9862
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 15198 7984 15254 7993
rect 15198 7919 15254 7928
rect 15212 7818 15240 7919
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 14830 7712 14886 7721
rect 14294 7644 14602 7653
rect 14830 7647 14886 7656
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 14200 7500 14320 7528
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14108 6458 14136 7346
rect 14188 6792 14240 6798
rect 14186 6760 14188 6769
rect 14240 6760 14242 6769
rect 14186 6695 14242 6704
rect 14292 6662 14320 7500
rect 14844 7002 14872 7647
rect 15120 7410 15148 7754
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15120 7002 15148 7346
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 4434 14136 6054
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5302 14228 5646
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14108 4406 14228 4434
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 13820 3062 13872 3068
rect 14002 3088 14058 3097
rect 13544 3052 13596 3058
rect 14002 3023 14058 3032
rect 13544 2994 13596 3000
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 13360 2032 13412 2038
rect 13360 1974 13412 1980
rect 13648 800 13676 2790
rect 13726 2680 13782 2689
rect 13726 2615 13782 2624
rect 13740 2446 13768 2615
rect 14108 2514 14136 3334
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 1970 14136 2246
rect 14200 2106 14228 4406
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 14660 2378 14688 6598
rect 14752 4826 14780 6598
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 14476 870 14596 898
rect 14476 800 14504 870
rect 3790 368 3846 377
rect 3790 303 3846 312
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 14568 762 14596 870
rect 14752 762 14780 2586
rect 14844 2310 14872 6666
rect 15016 6316 15068 6322
rect 15120 6304 15148 6938
rect 15396 6798 15424 8570
rect 15488 8498 15516 10066
rect 15672 9654 15700 13670
rect 16132 12714 16160 13738
rect 16518 13628 16826 13637
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16776 12850 16804 13398
rect 17052 13297 17080 14350
rect 17144 14006 17172 14855
rect 17498 14512 17554 14521
rect 17498 14447 17554 14456
rect 17512 14006 17540 14447
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17696 14113 17724 14350
rect 17682 14104 17738 14113
rect 17682 14039 17738 14048
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17696 13705 17724 13806
rect 17682 13696 17738 13705
rect 17604 13654 17682 13682
rect 17038 13288 17094 13297
rect 17038 13223 17094 13232
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16132 12170 16160 12650
rect 16316 12434 16344 12786
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16224 12406 16344 12434
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16028 12096 16080 12102
rect 16224 12073 16252 12406
rect 16304 12096 16356 12102
rect 16028 12038 16080 12044
rect 16210 12064 16266 12073
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11218 15792 11494
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15764 11121 15792 11154
rect 15750 11112 15806 11121
rect 15750 11047 15806 11056
rect 15856 10742 15884 11562
rect 15948 11218 15976 12038
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15936 11008 15988 11014
rect 15934 10976 15936 10985
rect 15988 10976 15990 10985
rect 15934 10911 15990 10920
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10198 15792 10406
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9722 15792 9862
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 8566 15608 9454
rect 15672 8634 15700 9590
rect 15750 9208 15806 9217
rect 15750 9143 15752 9152
rect 15804 9143 15806 9152
rect 15752 9114 15804 9120
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15580 8401 15608 8502
rect 15566 8392 15622 8401
rect 15566 8327 15622 8336
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15488 7410 15516 8026
rect 15672 7886 15700 8230
rect 15764 8090 15792 8774
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15068 6276 15148 6304
rect 15016 6258 15068 6264
rect 15120 5710 15148 6276
rect 15488 5914 15516 7346
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15672 6225 15700 7142
rect 15658 6216 15714 6225
rect 15658 6151 15714 6160
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 5522 15148 5646
rect 15212 5642 15332 5658
rect 15200 5636 15332 5642
rect 15252 5630 15332 5636
rect 15200 5578 15252 5584
rect 15120 5494 15240 5522
rect 15212 4826 15240 5494
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 15120 1034 15148 4490
rect 15212 4214 15240 4762
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 15212 3738 15240 4150
rect 15304 4078 15332 5630
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15198 1048 15254 1057
rect 15120 1006 15198 1034
rect 15198 983 15254 992
rect 15304 800 15332 3878
rect 15382 3496 15438 3505
rect 15382 3431 15384 3440
rect 15436 3431 15438 3440
rect 15384 3402 15436 3408
rect 15488 3346 15516 5510
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15580 4282 15608 4694
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15580 3466 15608 4218
rect 15672 4078 15700 5170
rect 15764 4622 15792 7142
rect 15856 6458 15884 10678
rect 16040 10538 16068 12038
rect 16304 12038 16356 12044
rect 16210 11999 16266 12008
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 10810 16160 11494
rect 16224 11150 16252 11630
rect 16316 11150 16344 12038
rect 16408 11665 16436 12582
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11694 16528 12106
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16488 11688 16540 11694
rect 16394 11656 16450 11665
rect 16488 11630 16540 11636
rect 16394 11591 16450 11600
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 11354 16436 11494
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 16868 11354 16896 11698
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16304 11144 16356 11150
rect 16580 11144 16632 11150
rect 16304 11086 16356 11092
rect 16408 11092 16580 11098
rect 16408 11086 16632 11092
rect 16762 11112 16818 11121
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16132 10282 16160 10746
rect 16040 10254 16160 10282
rect 15934 10024 15990 10033
rect 15934 9959 15990 9968
rect 15948 9217 15976 9959
rect 16040 9625 16068 10254
rect 16118 10024 16174 10033
rect 16118 9959 16174 9968
rect 16026 9616 16082 9625
rect 16026 9551 16082 9560
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15934 9208 15990 9217
rect 15934 9143 15990 9152
rect 16040 8974 16068 9454
rect 16132 9042 16160 9959
rect 16224 9489 16252 11086
rect 16316 9625 16344 11086
rect 16408 11070 16620 11086
rect 16672 11076 16724 11082
rect 16408 10033 16436 11070
rect 16762 11047 16818 11056
rect 16672 11018 16724 11024
rect 16684 10810 16712 11018
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16776 10674 16804 11047
rect 16854 10976 16910 10985
rect 16854 10911 16910 10920
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16394 10024 16450 10033
rect 16394 9959 16450 9968
rect 16486 9888 16542 9897
rect 16486 9823 16542 9832
rect 16500 9722 16528 9823
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16302 9616 16358 9625
rect 16302 9551 16358 9560
rect 16210 9480 16266 9489
rect 16210 9415 16266 9424
rect 16302 9208 16358 9217
rect 16302 9143 16358 9152
rect 16316 9042 16344 9143
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16132 8650 16160 8978
rect 16408 8974 16436 9658
rect 16868 9586 16896 10911
rect 16960 10849 16988 11494
rect 17052 11098 17080 12582
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17144 11898 17172 12038
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17236 11830 17264 13126
rect 17512 12918 17540 13194
rect 17604 12986 17632 13654
rect 17682 13631 17738 13640
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17684 13320 17736 13326
rect 17682 13288 17684 13297
rect 17736 13288 17738 13297
rect 17682 13223 17738 13232
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17500 12912 17552 12918
rect 17498 12880 17500 12889
rect 17552 12880 17554 12889
rect 17316 12844 17368 12850
rect 17498 12815 17554 12824
rect 17316 12786 17368 12792
rect 17512 12789 17540 12815
rect 17328 12288 17356 12786
rect 17684 12776 17736 12782
rect 17590 12744 17646 12753
rect 17684 12718 17736 12724
rect 17590 12679 17646 12688
rect 17604 12646 17632 12679
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17328 12260 17448 12288
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11218 17172 11630
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17052 11070 17356 11098
rect 17420 11082 17448 12260
rect 17512 11762 17540 12582
rect 17696 12481 17724 12718
rect 17682 12472 17738 12481
rect 17682 12407 17738 12416
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17500 11212 17552 11218
rect 17604 11200 17632 12242
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17788 12186 17816 13398
rect 17880 12442 17908 14350
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 17958 13424 18014 13433
rect 17958 13359 17960 13368
rect 18012 13359 18014 13368
rect 17960 13330 18012 13336
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17972 12374 18000 13330
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17960 12232 18012 12238
rect 17958 12200 17960 12209
rect 18012 12200 18014 12209
rect 17696 12073 17724 12174
rect 17788 12158 17908 12186
rect 17776 12096 17828 12102
rect 17682 12064 17738 12073
rect 17776 12038 17828 12044
rect 17682 11999 17738 12008
rect 17552 11172 17632 11200
rect 17500 11154 17552 11160
rect 17040 11008 17092 11014
rect 17038 10976 17040 10985
rect 17224 11008 17276 11014
rect 17092 10976 17094 10985
rect 17224 10950 17276 10956
rect 17038 10911 17094 10920
rect 16946 10840 17002 10849
rect 17236 10810 17264 10950
rect 16946 10775 17002 10784
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17328 10690 17356 11070
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17328 10662 17448 10690
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 16960 9761 16988 10542
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17052 10062 17080 10406
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17040 9920 17092 9926
rect 17038 9888 17040 9897
rect 17092 9888 17094 9897
rect 17038 9823 17094 9832
rect 16946 9752 17002 9761
rect 16946 9687 17002 9696
rect 16856 9580 16908 9586
rect 16908 9540 16988 9568
rect 16856 9522 16908 9528
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16960 9110 16988 9540
rect 16948 9104 17000 9110
rect 17000 9064 17080 9092
rect 16948 9046 17000 9052
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16396 8968 16448 8974
rect 16210 8936 16266 8945
rect 16396 8910 16448 8916
rect 16210 8871 16266 8880
rect 16224 8838 16252 8871
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16132 8622 16252 8650
rect 16684 8634 16712 8774
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15948 7818 15976 8298
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16040 7546 16068 7754
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15948 6730 15976 6938
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15672 3754 15700 4014
rect 15672 3738 15792 3754
rect 15672 3732 15804 3738
rect 15672 3726 15752 3732
rect 15752 3674 15804 3680
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15488 3318 15608 3346
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15488 2514 15516 3062
rect 15580 3058 15608 3318
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15580 2582 15608 2790
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15856 1873 15884 5510
rect 15948 5234 15976 5782
rect 16040 5681 16068 7278
rect 16132 6730 16160 7346
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16224 6662 16252 8622
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16776 8401 16804 8434
rect 16762 8392 16818 8401
rect 16396 8356 16448 8362
rect 16762 8327 16818 8336
rect 16396 8298 16448 8304
rect 16408 7834 16436 8298
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16762 7984 16818 7993
rect 16762 7919 16818 7928
rect 16316 7806 16436 7834
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16316 6322 16344 7806
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 6390 16436 7686
rect 16776 7546 16804 7919
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16776 7290 16804 7482
rect 16868 7449 16896 8978
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16854 7440 16910 7449
rect 16854 7375 16910 7384
rect 16776 7262 16896 7290
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16670 6896 16726 6905
rect 16670 6831 16726 6840
rect 16684 6798 16712 6831
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16868 6322 16896 7262
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16026 5672 16082 5681
rect 16026 5607 16082 5616
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16040 4554 16068 5607
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15842 1864 15898 1873
rect 15384 1828 15436 1834
rect 15842 1799 15898 1808
rect 15384 1770 15436 1776
rect 15396 1465 15424 1770
rect 15382 1456 15438 1465
rect 15382 1391 15438 1400
rect 14568 734 14780 762
rect 15290 0 15346 800
rect 15948 649 15976 4422
rect 16040 3194 16068 4490
rect 16132 4214 16160 5510
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 16224 4078 16252 5850
rect 16316 5370 16344 6258
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16868 5914 16896 6258
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16764 5840 16816 5846
rect 16578 5808 16634 5817
rect 16396 5772 16448 5778
rect 16764 5782 16816 5788
rect 16578 5743 16634 5752
rect 16396 5714 16448 5720
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4729 16344 4966
rect 16408 4758 16436 5714
rect 16592 5234 16620 5743
rect 16776 5574 16804 5782
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16776 5166 16804 5510
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16396 4752 16448 4758
rect 16302 4720 16358 4729
rect 16396 4694 16448 4700
rect 16302 4655 16358 4664
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16316 4026 16344 4422
rect 16408 4282 16436 4422
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16776 4214 16804 4762
rect 16868 4690 16896 5510
rect 16960 5302 16988 8910
rect 17052 8634 17080 9064
rect 17144 8634 17172 10542
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17144 7313 17172 7482
rect 17130 7304 17186 7313
rect 17130 7239 17186 7248
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 17052 6322 17080 6870
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 17052 5953 17080 6054
rect 17038 5944 17094 5953
rect 17038 5879 17094 5888
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 17038 5264 17094 5273
rect 17038 5199 17094 5208
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16316 3998 16436 4026
rect 16304 3936 16356 3942
rect 16118 3904 16174 3913
rect 16304 3878 16356 3884
rect 16118 3839 16174 3848
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16132 800 16160 3839
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 2650 16252 3470
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16316 2446 16344 3878
rect 16408 3058 16436 3998
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16868 3194 16896 4422
rect 16960 4282 16988 5102
rect 17052 4826 17080 5199
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17038 4312 17094 4321
rect 16948 4276 17000 4282
rect 17038 4247 17094 4256
rect 16948 4218 17000 4224
rect 17052 4010 17080 4247
rect 17040 4004 17092 4010
rect 17040 3946 17092 3952
rect 17144 3194 17172 4558
rect 17236 4146 17264 10406
rect 17420 10062 17448 10662
rect 17512 10606 17540 11154
rect 17684 11144 17736 11150
rect 17590 11112 17646 11121
rect 17684 11086 17736 11092
rect 17590 11047 17646 11056
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17604 10418 17632 11047
rect 17696 10849 17724 11086
rect 17682 10840 17738 10849
rect 17682 10775 17738 10784
rect 17788 10690 17816 12038
rect 17880 11778 17908 12158
rect 17958 12135 18014 12144
rect 17880 11750 18000 11778
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17972 11506 18000 11750
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18064 11665 18092 11698
rect 18050 11656 18106 11665
rect 18050 11591 18106 11600
rect 17880 11121 17908 11494
rect 17972 11478 18092 11506
rect 17960 11144 18012 11150
rect 17866 11112 17922 11121
rect 17960 11086 18012 11092
rect 17866 11047 17922 11056
rect 17972 10713 18000 11086
rect 18064 10810 18092 11478
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17512 10390 17632 10418
rect 17696 10662 17816 10690
rect 17958 10704 18014 10713
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17328 8090 17356 9590
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17328 7002 17356 7890
rect 17420 7886 17448 9386
rect 17512 8498 17540 10390
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17604 9042 17632 10134
rect 17696 9654 17724 10662
rect 18156 10674 18184 12582
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 17958 10639 18014 10648
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 18050 10568 18106 10577
rect 17880 10441 17908 10542
rect 18050 10503 18106 10512
rect 17866 10432 17922 10441
rect 17866 10367 17922 10376
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17682 9072 17738 9081
rect 17592 9036 17644 9042
rect 17682 9007 17738 9016
rect 17592 8978 17644 8984
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17498 8392 17554 8401
rect 17498 8327 17500 8336
rect 17552 8327 17554 8336
rect 17500 8298 17552 8304
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17512 7834 17540 8026
rect 17604 7954 17632 8978
rect 17696 8634 17724 9007
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17684 7880 17736 7886
rect 17512 7806 17632 7834
rect 17684 7822 17736 7828
rect 17500 7744 17552 7750
rect 17498 7712 17500 7721
rect 17552 7712 17554 7721
rect 17498 7647 17554 7656
rect 17604 7478 17632 7806
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17420 6440 17448 7210
rect 17604 6866 17632 7278
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17420 6412 17540 6440
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17328 5710 17356 6054
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17316 5704 17368 5710
rect 17420 5681 17448 5714
rect 17316 5646 17368 5652
rect 17406 5672 17462 5681
rect 17512 5642 17540 6412
rect 17604 5846 17632 6802
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17406 5607 17462 5616
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17328 5370 17356 5510
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17328 4690 17356 5102
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17328 4078 17356 4626
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17222 3904 17278 3913
rect 17222 3839 17278 3848
rect 17236 3738 17264 3839
rect 17420 3738 17448 4490
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17406 3632 17462 3641
rect 17406 3567 17462 3576
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2683 16826 2692
rect 16868 2514 16896 2790
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17420 2446 17448 3567
rect 17512 3040 17540 5238
rect 17696 4622 17724 7822
rect 17788 7041 17816 9862
rect 17880 9761 17908 10066
rect 18064 10062 18092 10503
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17866 9752 17922 9761
rect 17866 9687 17922 9696
rect 17972 9602 18000 9930
rect 17880 9574 18000 9602
rect 17880 9450 17908 9574
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17972 8906 18000 9454
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 7886 17908 8774
rect 18064 8673 18092 8910
rect 18050 8664 18106 8673
rect 18050 8599 18106 8608
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17868 7880 17920 7886
rect 17972 7857 18000 8434
rect 17868 7822 17920 7828
rect 17958 7848 18014 7857
rect 17958 7783 18014 7792
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17774 7032 17830 7041
rect 17774 6967 17830 6976
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17788 6118 17816 6802
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17590 4448 17646 4457
rect 17590 4383 17646 4392
rect 17604 4214 17632 4383
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17696 3602 17724 4558
rect 17788 3670 17816 6054
rect 17880 4690 17908 7686
rect 18064 7585 18092 7686
rect 18050 7576 18106 7585
rect 18050 7511 18106 7520
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6866 18092 7278
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17972 4010 18000 6734
rect 18050 6352 18106 6361
rect 18050 6287 18052 6296
rect 18104 6287 18106 6296
rect 18052 6258 18104 6264
rect 18156 5658 18184 10134
rect 18248 9382 18276 11494
rect 18340 10169 18368 13806
rect 18800 13190 18828 16400
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18432 11257 18460 11698
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18510 10976 18566 10985
rect 18510 10911 18566 10920
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18432 10441 18460 10474
rect 18418 10432 18474 10441
rect 18418 10367 18474 10376
rect 18326 10160 18382 10169
rect 18326 10095 18382 10104
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18432 9722 18460 10066
rect 18524 9994 18552 10911
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 7750 18276 8910
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18340 7970 18368 8842
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18418 8392 18474 8401
rect 18418 8327 18474 8336
rect 18432 8090 18460 8327
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18524 7993 18552 8774
rect 18510 7984 18566 7993
rect 18340 7942 18460 7970
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18432 7834 18460 7942
rect 18510 7919 18566 7928
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18340 7546 18368 7822
rect 18432 7806 18552 7834
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18418 7168 18474 7177
rect 18418 7103 18474 7112
rect 18432 7002 18460 7103
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18418 6760 18474 6769
rect 18248 6458 18276 6734
rect 18328 6724 18380 6730
rect 18418 6695 18474 6704
rect 18328 6666 18380 6672
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18248 6225 18276 6258
rect 18234 6216 18290 6225
rect 18234 6151 18290 6160
rect 18064 5630 18184 5658
rect 18064 4622 18092 5630
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18156 4826 18184 5510
rect 18248 5370 18276 5510
rect 18340 5370 18368 6666
rect 18432 6662 18460 6695
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18432 6361 18460 6394
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18524 6066 18552 7806
rect 18616 6934 18644 9386
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18524 6038 18644 6066
rect 18418 5536 18474 5545
rect 18418 5471 18474 5480
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17788 3398 17816 3606
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17592 3052 17644 3058
rect 17512 3012 17592 3040
rect 17592 2994 17644 3000
rect 17788 2990 17816 3334
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 17972 2922 18000 3402
rect 18050 3088 18106 3097
rect 18050 3023 18106 3032
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17498 2680 17554 2689
rect 17498 2615 17554 2624
rect 17774 2680 17830 2689
rect 18064 2650 18092 3023
rect 18248 2774 18276 4966
rect 18340 3738 18368 5034
rect 18432 4826 18460 5471
rect 18616 5234 18644 6038
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18510 5128 18566 5137
rect 18510 5063 18566 5072
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18524 4282 18552 5063
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18616 4162 18644 5170
rect 18524 4134 18644 4162
rect 18708 4146 18736 11562
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18696 4140 18748 4146
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18418 3496 18474 3505
rect 18418 3431 18474 3440
rect 18156 2746 18276 2774
rect 17774 2615 17776 2624
rect 17512 2446 17540 2615
rect 17828 2615 17830 2624
rect 18052 2644 18104 2650
rect 17776 2586 17828 2592
rect 18052 2586 18104 2592
rect 18156 2446 18184 2746
rect 18432 2650 18460 3431
rect 18524 3194 18552 4134
rect 18696 4082 18748 4088
rect 18602 4040 18658 4049
rect 18602 3975 18658 3984
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 16948 2304 17000 2310
rect 16946 2272 16948 2281
rect 17776 2304 17828 2310
rect 17000 2272 17002 2281
rect 17776 2246 17828 2252
rect 16946 2207 17002 2216
rect 16948 2032 17000 2038
rect 16948 1974 17000 1980
rect 16960 800 16988 1974
rect 17788 800 17816 2246
rect 17880 2106 17908 2382
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 18616 800 18644 3975
rect 18800 3602 18828 8298
rect 18892 4078 18920 8366
rect 18984 5166 19012 11222
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18984 3534 19012 5102
rect 19076 4690 19104 7278
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 15934 640 15990 649
rect 15934 575 15990 584
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
<< via2 >>
rect 4434 16632 4490 16688
rect 2962 15408 3018 15464
rect 1490 11328 1546 11384
rect 1490 10512 1546 10568
rect 1306 8336 1362 8392
rect 2226 14184 2282 14240
rect 2226 13776 2282 13832
rect 2778 14612 2834 14648
rect 2778 14592 2780 14612
rect 2780 14592 2832 14612
rect 2832 14592 2834 14612
rect 3054 15000 3110 15056
rect 3698 16224 3754 16280
rect 3606 15816 3662 15872
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 2870 13812 2872 13832
rect 2872 13812 2924 13832
rect 2924 13812 2926 13832
rect 3330 13912 3386 13968
rect 2870 13776 2926 13812
rect 2778 13368 2834 13424
rect 1950 12280 2006 12336
rect 1674 9968 1730 10024
rect 1490 9832 1546 9888
rect 1490 8880 1546 8936
rect 1766 8780 1768 8800
rect 1768 8780 1820 8800
rect 1820 8780 1822 8800
rect 1766 8744 1822 8780
rect 1766 8608 1822 8664
rect 1490 8084 1546 8120
rect 1490 8064 1492 8084
rect 1492 8064 1544 8084
rect 1544 8064 1546 8084
rect 1490 7268 1546 7304
rect 1490 7248 1492 7268
rect 1492 7248 1544 7268
rect 1544 7248 1546 7268
rect 1490 6876 1492 6896
rect 1492 6876 1544 6896
rect 1544 6876 1546 6896
rect 1490 6840 1546 6876
rect 2042 11736 2098 11792
rect 2226 12552 2282 12608
rect 2226 12180 2228 12200
rect 2228 12180 2280 12200
rect 2280 12180 2282 12200
rect 2226 12144 2282 12180
rect 1950 11056 2006 11112
rect 2042 7928 2098 7984
rect 2226 10920 2282 10976
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 2870 12960 2926 13016
rect 3146 13268 3148 13288
rect 3148 13268 3200 13288
rect 3200 13268 3202 13288
rect 3146 13232 3202 13268
rect 2962 12824 3018 12880
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 2962 12416 3018 12472
rect 2778 11736 2834 11792
rect 2502 11192 2558 11248
rect 2410 10920 2466 10976
rect 2226 9696 2282 9752
rect 2870 9696 2926 9752
rect 3514 12144 3570 12200
rect 3054 11736 3110 11792
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 3054 10648 3110 10704
rect 3974 13776 4030 13832
rect 3790 13504 3846 13560
rect 3698 13368 3754 13424
rect 4066 13368 4122 13424
rect 4158 13252 4214 13288
rect 4158 13232 4160 13252
rect 4160 13232 4212 13252
rect 4212 13232 4214 13252
rect 3606 10648 3662 10704
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3054 10104 3110 10160
rect 3606 10376 3662 10432
rect 2410 8880 2466 8936
rect 2318 8608 2374 8664
rect 1858 7692 1860 7712
rect 1860 7692 1912 7712
rect 1912 7692 1914 7712
rect 1858 7656 1914 7692
rect 1858 6432 1914 6488
rect 2226 7420 2228 7440
rect 2228 7420 2280 7440
rect 2280 7420 2282 7440
rect 2226 7384 2282 7420
rect 3054 9560 3110 9616
rect 3514 9832 3570 9888
rect 3790 11348 3846 11384
rect 3790 11328 3792 11348
rect 3792 11328 3844 11348
rect 3844 11328 3846 11348
rect 4894 14320 4950 14376
rect 4342 12688 4398 12744
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 16302 16496 16358 16552
rect 16026 16088 16082 16144
rect 7378 13912 7434 13968
rect 5722 13640 5778 13696
rect 3974 10804 4030 10840
rect 3974 10784 3976 10804
rect 3976 10784 4028 10804
rect 4028 10784 4030 10804
rect 3974 9696 4030 9752
rect 2502 6840 2558 6896
rect 1490 6060 1492 6080
rect 1492 6060 1544 6080
rect 1544 6060 1546 6080
rect 1490 6024 1546 6060
rect 1582 5616 1638 5672
rect 1122 3304 1178 3360
rect 1674 5480 1730 5536
rect 1490 5208 1546 5264
rect 1490 4800 1546 4856
rect 1490 4428 1492 4448
rect 1492 4428 1544 4448
rect 1544 4428 1546 4448
rect 1490 4392 1546 4428
rect 1490 4004 1546 4040
rect 1490 3984 1492 4004
rect 1492 3984 1544 4004
rect 1544 3984 1546 4004
rect 1674 3984 1730 4040
rect 1490 3168 1546 3224
rect 2226 6160 2282 6216
rect 2134 5208 2190 5264
rect 1950 4664 2006 4720
rect 1858 3576 1914 3632
rect 2042 3848 2098 3904
rect 1582 2760 1638 2816
rect 1858 2352 1914 2408
rect 2042 2760 2098 2816
rect 1950 1128 2006 1184
rect 2870 9288 2926 9344
rect 3606 9424 3662 9480
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3330 9016 3386 9072
rect 2962 8472 3018 8528
rect 3422 8372 3424 8392
rect 3424 8372 3476 8392
rect 3476 8372 3478 8392
rect 3422 8336 3478 8372
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3146 7248 3202 7304
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3330 6704 3386 6760
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 3146 5752 3202 5808
rect 3054 5616 3110 5672
rect 2594 3440 2650 3496
rect 2226 1944 2282 2000
rect 3422 5480 3478 5536
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 3054 3984 3110 4040
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 2686 1536 2742 1592
rect 3606 7928 3662 7984
rect 3790 8744 3846 8800
rect 3882 8472 3938 8528
rect 3606 6024 3662 6080
rect 3422 3052 3478 3088
rect 3422 3032 3424 3052
rect 3424 3032 3476 3052
rect 3476 3032 3478 3052
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 1674 720 1730 776
rect 4158 11328 4214 11384
rect 4250 9988 4306 10024
rect 4250 9968 4252 9988
rect 4252 9968 4304 9988
rect 4304 9968 4306 9988
rect 4894 13368 4950 13424
rect 5814 13368 5870 13424
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 5998 12824 6054 12880
rect 4986 12688 5042 12744
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 4986 11600 5042 11656
rect 4986 11056 5042 11112
rect 4986 10956 4988 10976
rect 4988 10956 5040 10976
rect 5040 10956 5042 10976
rect 4986 10920 5042 10956
rect 4986 10804 5042 10840
rect 4986 10784 4988 10804
rect 4988 10784 5040 10804
rect 5040 10784 5042 10804
rect 5814 11328 5870 11384
rect 4986 10512 5042 10568
rect 4618 10376 4674 10432
rect 4986 10240 5042 10296
rect 4158 9288 4214 9344
rect 4158 8608 4214 8664
rect 4526 9460 4528 9480
rect 4528 9460 4580 9480
rect 4580 9460 4582 9480
rect 4526 9424 4582 9460
rect 4894 9832 4950 9888
rect 5170 10376 5226 10432
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5814 10804 5870 10840
rect 5814 10784 5816 10804
rect 5816 10784 5868 10804
rect 5868 10784 5870 10804
rect 5262 10240 5318 10296
rect 5446 9968 5502 10024
rect 5722 9968 5778 10024
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 6826 13524 6882 13560
rect 6826 13504 6828 13524
rect 6828 13504 6880 13524
rect 6880 13504 6882 13524
rect 6366 12824 6422 12880
rect 6550 12144 6606 12200
rect 4158 7964 4160 7984
rect 4160 7964 4212 7984
rect 4212 7964 4214 7984
rect 4158 7928 4214 7964
rect 4066 7384 4122 7440
rect 4158 6724 4214 6760
rect 4158 6704 4160 6724
rect 4160 6704 4212 6724
rect 4212 6704 4214 6724
rect 4342 7520 4398 7576
rect 4434 7384 4490 7440
rect 4342 6296 4398 6352
rect 4342 5888 4398 5944
rect 4158 5616 4214 5672
rect 3882 2644 3938 2680
rect 3882 2624 3884 2644
rect 3884 2624 3936 2644
rect 3936 2624 3938 2644
rect 4802 6024 4858 6080
rect 4710 5752 4766 5808
rect 4342 3340 4344 3360
rect 4344 3340 4396 3360
rect 4396 3340 4398 3360
rect 4342 3304 4398 3340
rect 4342 2896 4398 2952
rect 5998 9288 6054 9344
rect 5906 9152 5962 9208
rect 5630 9036 5686 9072
rect 5630 9016 5632 9036
rect 5632 9016 5684 9036
rect 5684 9016 5686 9036
rect 5814 8916 5816 8936
rect 5816 8916 5868 8936
rect 5868 8916 5870 8936
rect 5814 8880 5870 8916
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5078 7792 5134 7848
rect 5722 7828 5724 7848
rect 5724 7828 5776 7848
rect 5776 7828 5778 7848
rect 5722 7792 5778 7828
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5538 7404 5594 7440
rect 5538 7384 5540 7404
rect 5540 7384 5592 7404
rect 5592 7384 5594 7404
rect 5722 6840 5778 6896
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5170 5888 5226 5944
rect 5814 6160 5870 6216
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 4802 2760 4858 2816
rect 6366 10376 6422 10432
rect 6366 9288 6422 9344
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 6826 11092 6828 11112
rect 6828 11092 6880 11112
rect 6880 11092 6882 11112
rect 6826 11056 6882 11092
rect 6642 9696 6698 9752
rect 6274 9016 6330 9072
rect 6274 4664 6330 4720
rect 6090 3052 6146 3088
rect 6090 3032 6092 3052
rect 6092 3032 6144 3052
rect 6144 3032 6146 3052
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 6550 8200 6606 8256
rect 6826 9832 6882 9888
rect 7194 11056 7250 11112
rect 6734 5616 6790 5672
rect 6734 5208 6790 5264
rect 7102 5072 7158 5128
rect 6918 4120 6974 4176
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 7470 9832 7526 9888
rect 7930 9696 7986 9752
rect 7838 9560 7894 9616
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 7378 6024 7434 6080
rect 8022 8336 8078 8392
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 8666 9560 8722 9616
rect 8574 9016 8630 9072
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 9586 13232 9642 13288
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9402 12008 9458 12064
rect 9218 11636 9220 11656
rect 9220 11636 9272 11656
rect 9272 11636 9274 11656
rect 9218 11600 9274 11636
rect 10506 13776 10562 13832
rect 9678 12280 9734 12336
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9402 11600 9458 11656
rect 9310 11500 9312 11520
rect 9312 11500 9364 11520
rect 9364 11500 9366 11520
rect 9310 11464 9366 11500
rect 9218 11056 9274 11112
rect 9034 10784 9090 10840
rect 10230 11192 10286 11248
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9494 8472 9550 8528
rect 9310 7928 9366 7984
rect 9402 3576 9458 3632
rect 8114 2932 8116 2952
rect 8116 2932 8168 2952
rect 8168 2932 8170 2952
rect 8114 2896 8170 2932
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10230 9424 10286 9480
rect 9770 9016 9826 9072
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10230 7928 10286 7984
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10414 12008 10470 12064
rect 10414 11228 10416 11248
rect 10416 11228 10468 11248
rect 10468 11228 10470 11248
rect 10414 11192 10470 11228
rect 10782 11600 10838 11656
rect 10138 4664 10194 4720
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10598 5616 10654 5672
rect 10598 4120 10654 4176
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9402 2488 9458 2544
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 11794 12688 11850 12744
rect 10966 4528 11022 4584
rect 11334 10668 11390 10704
rect 11334 10648 11336 10668
rect 11336 10648 11388 10668
rect 11388 10648 11390 10668
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 12530 12436 12586 12472
rect 12530 12416 12532 12436
rect 12532 12416 12584 12436
rect 12584 12416 12586 12436
rect 11794 11736 11850 11792
rect 11702 10648 11758 10704
rect 11426 10104 11482 10160
rect 11334 9036 11390 9072
rect 11334 9016 11336 9036
rect 11336 9016 11388 9036
rect 11388 9016 11390 9036
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 11702 9968 11758 10024
rect 11886 10004 11888 10024
rect 11888 10004 11940 10024
rect 11940 10004 11942 10024
rect 11886 9968 11942 10004
rect 11794 9016 11850 9072
rect 11150 5208 11206 5264
rect 11610 8336 11666 8392
rect 11702 7248 11758 7304
rect 11702 6568 11758 6624
rect 11150 3984 11206 4040
rect 11242 3440 11298 3496
rect 11702 5616 11758 5672
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12438 10104 12494 10160
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12162 6704 12218 6760
rect 12438 6704 12494 6760
rect 12438 6568 12494 6624
rect 12254 6452 12310 6488
rect 12254 6432 12256 6452
rect 12256 6432 12308 6452
rect 12308 6432 12310 6452
rect 12162 6296 12218 6352
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 12254 5772 12310 5808
rect 12254 5752 12256 5772
rect 12256 5752 12308 5772
rect 12308 5752 12310 5772
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 12346 3984 12402 4040
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 13542 13812 13544 13832
rect 13544 13812 13596 13832
rect 13596 13812 13598 13832
rect 13542 13776 13598 13812
rect 13450 13232 13506 13288
rect 12990 7792 13046 7848
rect 12898 7384 12954 7440
rect 12990 6860 13046 6896
rect 12990 6840 12992 6860
rect 12992 6840 13044 6860
rect 13044 6840 13046 6860
rect 12806 6316 12862 6352
rect 12990 6432 13046 6488
rect 12806 6296 12808 6316
rect 12808 6296 12860 6316
rect 12860 6296 12862 6316
rect 13450 12860 13452 12880
rect 13452 12860 13504 12880
rect 13504 12860 13506 12880
rect 13450 12824 13506 12860
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 15474 14492 15476 14512
rect 15476 14492 15528 14512
rect 15528 14492 15530 14512
rect 15474 14456 15530 14492
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14094 12960 14150 13016
rect 14554 12416 14610 12472
rect 13266 9424 13322 9480
rect 16210 15680 16266 15736
rect 16394 15272 16450 15328
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 17130 14864 17186 14920
rect 16670 14320 16726 14376
rect 15474 13776 15530 13832
rect 16854 13796 16910 13832
rect 16854 13776 16856 13796
rect 16856 13776 16908 13796
rect 16908 13776 16910 13796
rect 15106 12416 15162 12472
rect 13818 12144 13874 12200
rect 13818 11872 13874 11928
rect 13450 9152 13506 9208
rect 13358 8472 13414 8528
rect 13634 8608 13690 8664
rect 13634 7828 13636 7848
rect 13636 7828 13688 7848
rect 13688 7828 13690 7848
rect 13634 7792 13690 7828
rect 13634 7520 13690 7576
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 14554 11192 14610 11248
rect 14094 11056 14150 11112
rect 14002 9696 14058 9752
rect 13542 7284 13544 7304
rect 13544 7284 13596 7304
rect 13596 7284 13598 7304
rect 13542 7248 13598 7284
rect 13634 6704 13690 6760
rect 12622 2896 12678 2952
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 13726 6568 13782 6624
rect 14002 8064 14058 8120
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14738 10784 14794 10840
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 14738 9696 14794 9752
rect 14370 9288 14426 9344
rect 14186 9152 14242 9208
rect 14462 9152 14518 9208
rect 15014 12280 15070 12336
rect 14830 9288 14886 9344
rect 14830 9036 14886 9072
rect 14830 9016 14832 9036
rect 14832 9016 14884 9036
rect 14884 9016 14886 9036
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14738 8608 14794 8664
rect 15566 10240 15622 10296
rect 15290 9832 15346 9888
rect 15198 8744 15254 8800
rect 15198 7928 15254 7984
rect 14830 7656 14886 7712
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14186 6740 14188 6760
rect 14188 6740 14240 6760
rect 14240 6740 14242 6760
rect 14186 6704 14242 6740
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14002 3032 14058 3088
rect 13726 2624 13782 2680
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 3790 312 3846 368
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 17498 14456 17554 14512
rect 17682 14048 17738 14104
rect 17038 13232 17094 13288
rect 15750 11056 15806 11112
rect 15934 10956 15936 10976
rect 15936 10956 15988 10976
rect 15988 10956 15990 10976
rect 15934 10920 15990 10956
rect 15750 9172 15806 9208
rect 15750 9152 15752 9172
rect 15752 9152 15804 9172
rect 15804 9152 15806 9172
rect 15566 8336 15622 8392
rect 15658 6160 15714 6216
rect 15198 992 15254 1048
rect 15382 3460 15438 3496
rect 15382 3440 15384 3460
rect 15384 3440 15436 3460
rect 15436 3440 15438 3460
rect 16210 12008 16266 12064
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16394 11600 16450 11656
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 15934 9968 15990 10024
rect 16118 9968 16174 10024
rect 16026 9560 16082 9616
rect 15934 9152 15990 9208
rect 16762 11056 16818 11112
rect 16854 10920 16910 10976
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16394 9968 16450 10024
rect 16486 9832 16542 9888
rect 16302 9560 16358 9616
rect 16210 9424 16266 9480
rect 16302 9152 16358 9208
rect 17682 13640 17738 13696
rect 17682 13268 17684 13288
rect 17684 13268 17736 13288
rect 17736 13268 17738 13288
rect 17682 13232 17738 13268
rect 17498 12860 17500 12880
rect 17500 12860 17552 12880
rect 17552 12860 17554 12880
rect 17498 12824 17554 12860
rect 17590 12688 17646 12744
rect 17682 12416 17738 12472
rect 17958 13388 18014 13424
rect 17958 13368 17960 13388
rect 17960 13368 18012 13388
rect 18012 13368 18014 13388
rect 17682 12008 17738 12064
rect 17038 10956 17040 10976
rect 17040 10956 17092 10976
rect 17092 10956 17094 10976
rect 17038 10920 17094 10956
rect 16946 10784 17002 10840
rect 17038 9868 17040 9888
rect 17040 9868 17092 9888
rect 17092 9868 17094 9888
rect 17038 9832 17094 9868
rect 16946 9696 17002 9752
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16210 8880 16266 8936
rect 16762 8336 16818 8392
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16762 7928 16818 7984
rect 16854 7384 16910 7440
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16670 6840 16726 6896
rect 16026 5616 16082 5672
rect 15842 1808 15898 1864
rect 15382 1400 15438 1456
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16578 5752 16634 5808
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16302 4664 16358 4720
rect 17130 7248 17186 7304
rect 17038 5888 17094 5944
rect 17038 5208 17094 5264
rect 16118 3848 16174 3904
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 17038 4256 17094 4312
rect 17590 11056 17646 11112
rect 17682 10784 17738 10840
rect 17958 12180 17960 12200
rect 17960 12180 18012 12200
rect 18012 12180 18014 12200
rect 17958 12144 18014 12180
rect 18050 11600 18106 11656
rect 17866 11056 17922 11112
rect 17958 10648 18014 10704
rect 18050 10512 18106 10568
rect 17866 10376 17922 10432
rect 17682 9016 17738 9072
rect 17498 8356 17554 8392
rect 17498 8336 17500 8356
rect 17500 8336 17552 8356
rect 17552 8336 17554 8356
rect 17498 7692 17500 7712
rect 17500 7692 17552 7712
rect 17552 7692 17554 7712
rect 17498 7656 17554 7692
rect 17406 5616 17462 5672
rect 17222 3848 17278 3904
rect 17406 3576 17462 3632
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 17866 9696 17922 9752
rect 18050 8608 18106 8664
rect 17958 7792 18014 7848
rect 17774 6976 17830 7032
rect 17590 4392 17646 4448
rect 18050 7520 18106 7576
rect 18050 6316 18106 6352
rect 18050 6296 18052 6316
rect 18052 6296 18104 6316
rect 18104 6296 18106 6316
rect 18418 11192 18474 11248
rect 18510 10920 18566 10976
rect 18418 10376 18474 10432
rect 18326 10104 18382 10160
rect 18418 8336 18474 8392
rect 18510 7928 18566 7984
rect 18418 7112 18474 7168
rect 18418 6704 18474 6760
rect 18234 6160 18290 6216
rect 18418 6296 18474 6352
rect 18418 5480 18474 5536
rect 18050 3032 18106 3088
rect 17498 2624 17554 2680
rect 17774 2644 17830 2680
rect 18510 5072 18566 5128
rect 18418 3440 18474 3496
rect 17774 2624 17776 2644
rect 17776 2624 17828 2644
rect 17828 2624 17830 2644
rect 18602 3984 18658 4040
rect 16946 2252 16948 2272
rect 16948 2252 17000 2272
rect 17000 2252 17002 2272
rect 16946 2216 17002 2252
rect 15934 584 15990 640
<< metal3 >>
rect 0 16690 800 16720
rect 4429 16690 4495 16693
rect 0 16688 4495 16690
rect 0 16632 4434 16688
rect 4490 16632 4495 16688
rect 0 16630 4495 16632
rect 0 16600 800 16630
rect 4429 16627 4495 16630
rect 16297 16554 16363 16557
rect 19200 16554 20000 16584
rect 16297 16552 20000 16554
rect 16297 16496 16302 16552
rect 16358 16496 20000 16552
rect 16297 16494 20000 16496
rect 16297 16491 16363 16494
rect 19200 16464 20000 16494
rect 0 16282 800 16312
rect 3693 16282 3759 16285
rect 0 16280 3759 16282
rect 0 16224 3698 16280
rect 3754 16224 3759 16280
rect 0 16222 3759 16224
rect 0 16192 800 16222
rect 3693 16219 3759 16222
rect 16021 16146 16087 16149
rect 19200 16146 20000 16176
rect 16021 16144 20000 16146
rect 16021 16088 16026 16144
rect 16082 16088 20000 16144
rect 16021 16086 20000 16088
rect 16021 16083 16087 16086
rect 19200 16056 20000 16086
rect 0 15874 800 15904
rect 3601 15874 3667 15877
rect 0 15872 3667 15874
rect 0 15816 3606 15872
rect 3662 15816 3667 15872
rect 0 15814 3667 15816
rect 0 15784 800 15814
rect 3601 15811 3667 15814
rect 16205 15738 16271 15741
rect 19200 15738 20000 15768
rect 16205 15736 20000 15738
rect 16205 15680 16210 15736
rect 16266 15680 20000 15736
rect 16205 15678 20000 15680
rect 16205 15675 16271 15678
rect 19200 15648 20000 15678
rect 0 15466 800 15496
rect 2957 15466 3023 15469
rect 0 15464 3023 15466
rect 0 15408 2962 15464
rect 3018 15408 3023 15464
rect 0 15406 3023 15408
rect 0 15376 800 15406
rect 2957 15403 3023 15406
rect 16389 15330 16455 15333
rect 19200 15330 20000 15360
rect 16389 15328 20000 15330
rect 16389 15272 16394 15328
rect 16450 15272 20000 15328
rect 16389 15270 20000 15272
rect 16389 15267 16455 15270
rect 19200 15240 20000 15270
rect 0 15058 800 15088
rect 3049 15058 3115 15061
rect 0 15056 3115 15058
rect 0 15000 3054 15056
rect 3110 15000 3115 15056
rect 0 14998 3115 15000
rect 0 14968 800 14998
rect 3049 14995 3115 14998
rect 17125 14922 17191 14925
rect 19200 14922 20000 14952
rect 17125 14920 20000 14922
rect 17125 14864 17130 14920
rect 17186 14864 20000 14920
rect 17125 14862 20000 14864
rect 17125 14859 17191 14862
rect 19200 14832 20000 14862
rect 3170 14720 3486 14721
rect 0 14650 800 14680
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 2773 14650 2839 14653
rect 0 14648 2839 14650
rect 0 14592 2778 14648
rect 2834 14592 2839 14648
rect 0 14590 2839 14592
rect 0 14560 800 14590
rect 2773 14587 2839 14590
rect 15469 14514 15535 14517
rect 17493 14514 17559 14517
rect 19200 14514 20000 14544
rect 15469 14512 20000 14514
rect 15469 14456 15474 14512
rect 15530 14456 17498 14512
rect 17554 14456 20000 14512
rect 15469 14454 20000 14456
rect 15469 14451 15535 14454
rect 17493 14451 17559 14454
rect 19200 14424 20000 14454
rect 4889 14378 4955 14381
rect 16665 14378 16731 14381
rect 4889 14376 16731 14378
rect 4889 14320 4894 14376
rect 4950 14320 16670 14376
rect 16726 14320 16731 14376
rect 4889 14318 16731 14320
rect 4889 14315 4955 14318
rect 16665 14315 16731 14318
rect 0 14242 800 14272
rect 2221 14242 2287 14245
rect 0 14240 2287 14242
rect 0 14184 2226 14240
rect 2282 14184 2287 14240
rect 0 14182 2287 14184
rect 0 14152 800 14182
rect 2221 14179 2287 14182
rect 5394 14176 5710 14177
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 14290 14111 14606 14112
rect 17677 14106 17743 14109
rect 19200 14106 20000 14136
rect 17677 14104 20000 14106
rect 17677 14048 17682 14104
rect 17738 14048 20000 14104
rect 17677 14046 20000 14048
rect 17677 14043 17743 14046
rect 19200 14016 20000 14046
rect 3325 13970 3391 13973
rect 3550 13970 3556 13972
rect 3325 13968 3556 13970
rect 3325 13912 3330 13968
rect 3386 13912 3556 13968
rect 3325 13910 3556 13912
rect 3325 13907 3391 13910
rect 3550 13908 3556 13910
rect 3620 13970 3626 13972
rect 7373 13970 7439 13973
rect 3620 13968 7439 13970
rect 3620 13912 7378 13968
rect 7434 13912 7439 13968
rect 3620 13910 7439 13912
rect 3620 13908 3626 13910
rect 7373 13907 7439 13910
rect 0 13834 800 13864
rect 2221 13834 2287 13837
rect 0 13832 2287 13834
rect 0 13776 2226 13832
rect 2282 13776 2287 13832
rect 0 13774 2287 13776
rect 0 13744 800 13774
rect 2221 13771 2287 13774
rect 2865 13834 2931 13837
rect 3969 13834 4035 13837
rect 10501 13834 10567 13837
rect 13537 13836 13603 13837
rect 13486 13834 13492 13836
rect 2865 13832 3802 13834
rect 2865 13776 2870 13832
rect 2926 13776 3802 13832
rect 2865 13774 3802 13776
rect 2865 13771 2931 13774
rect 3742 13698 3802 13774
rect 3969 13832 10567 13834
rect 3969 13776 3974 13832
rect 4030 13776 10506 13832
rect 10562 13776 10567 13832
rect 3969 13774 10567 13776
rect 13446 13774 13492 13834
rect 13556 13832 13603 13836
rect 13598 13776 13603 13832
rect 3969 13771 4035 13774
rect 10501 13771 10567 13774
rect 13486 13772 13492 13774
rect 13556 13772 13603 13776
rect 13670 13772 13676 13836
rect 13740 13834 13746 13836
rect 15469 13834 15535 13837
rect 13740 13832 15535 13834
rect 13740 13776 15474 13832
rect 15530 13776 15535 13832
rect 13740 13774 15535 13776
rect 13740 13772 13746 13774
rect 13537 13771 13603 13772
rect 15469 13771 15535 13774
rect 16849 13834 16915 13837
rect 17534 13834 17540 13836
rect 16849 13832 17540 13834
rect 16849 13776 16854 13832
rect 16910 13776 17540 13832
rect 16849 13774 17540 13776
rect 16849 13771 16915 13774
rect 17534 13772 17540 13774
rect 17604 13772 17610 13836
rect 5717 13698 5783 13701
rect 3742 13696 5783 13698
rect 3742 13640 5722 13696
rect 5778 13640 5783 13696
rect 3742 13638 5783 13640
rect 5717 13635 5783 13638
rect 17677 13698 17743 13701
rect 19200 13698 20000 13728
rect 17677 13696 20000 13698
rect 17677 13640 17682 13696
rect 17738 13640 20000 13696
rect 17677 13638 20000 13640
rect 17677 13635 17743 13638
rect 3170 13632 3486 13633
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 19200 13608 20000 13638
rect 16514 13567 16830 13568
rect 3785 13564 3851 13565
rect 3734 13500 3740 13564
rect 3804 13562 3851 13564
rect 6821 13562 6887 13565
rect 3804 13560 6887 13562
rect 3846 13504 6826 13560
rect 6882 13504 6887 13560
rect 3804 13502 6887 13504
rect 3804 13500 3851 13502
rect 3785 13499 3851 13500
rect 6821 13499 6887 13502
rect 0 13426 800 13456
rect 2773 13426 2839 13429
rect 0 13424 2839 13426
rect 0 13368 2778 13424
rect 2834 13368 2839 13424
rect 0 13366 2839 13368
rect 0 13336 800 13366
rect 2773 13363 2839 13366
rect 3693 13426 3759 13429
rect 4061 13426 4127 13429
rect 3693 13424 4127 13426
rect 3693 13368 3698 13424
rect 3754 13368 4066 13424
rect 4122 13368 4127 13424
rect 3693 13366 4127 13368
rect 3693 13363 3759 13366
rect 4061 13363 4127 13366
rect 4889 13426 4955 13429
rect 5809 13426 5875 13429
rect 17953 13426 18019 13429
rect 4889 13424 18019 13426
rect 4889 13368 4894 13424
rect 4950 13368 5814 13424
rect 5870 13368 17958 13424
rect 18014 13368 18019 13424
rect 4889 13366 18019 13368
rect 4889 13363 4955 13366
rect 5809 13363 5875 13366
rect 17953 13363 18019 13366
rect 3141 13290 3207 13293
rect 4153 13290 4219 13293
rect 9581 13290 9647 13293
rect 3141 13288 9647 13290
rect 3141 13232 3146 13288
rect 3202 13232 4158 13288
rect 4214 13232 9586 13288
rect 9642 13232 9647 13288
rect 3141 13230 9647 13232
rect 3141 13227 3207 13230
rect 4153 13227 4219 13230
rect 9581 13227 9647 13230
rect 13445 13290 13511 13293
rect 17033 13290 17099 13293
rect 13445 13288 17099 13290
rect 13445 13232 13450 13288
rect 13506 13232 17038 13288
rect 17094 13232 17099 13288
rect 13445 13230 17099 13232
rect 13445 13227 13511 13230
rect 17033 13227 17099 13230
rect 17677 13290 17743 13293
rect 19200 13290 20000 13320
rect 17677 13288 20000 13290
rect 17677 13232 17682 13288
rect 17738 13232 20000 13288
rect 17677 13230 20000 13232
rect 17677 13227 17743 13230
rect 19200 13200 20000 13230
rect 5394 13088 5710 13089
rect 0 13018 800 13048
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 14290 13023 14606 13024
rect 2865 13018 2931 13021
rect 14089 13018 14155 13021
rect 0 13016 2931 13018
rect 0 12960 2870 13016
rect 2926 12960 2931 13016
rect 0 12958 2931 12960
rect 0 12928 800 12958
rect 2865 12955 2931 12958
rect 10320 13016 14155 13018
rect 10320 12960 14094 13016
rect 14150 12960 14155 13016
rect 10320 12958 14155 12960
rect 2957 12882 3023 12885
rect 3918 12882 3924 12884
rect 2957 12880 3924 12882
rect 2957 12824 2962 12880
rect 3018 12824 3924 12880
rect 2957 12822 3924 12824
rect 2957 12819 3023 12822
rect 3918 12820 3924 12822
rect 3988 12882 3994 12884
rect 5993 12882 6059 12885
rect 6361 12884 6427 12885
rect 6310 12882 6316 12884
rect 3988 12880 6059 12882
rect 3988 12824 5998 12880
rect 6054 12824 6059 12880
rect 3988 12822 6059 12824
rect 6234 12822 6316 12882
rect 6380 12882 6427 12884
rect 10320 12882 10380 12958
rect 14089 12955 14155 12958
rect 13445 12882 13511 12885
rect 6380 12880 10380 12882
rect 6422 12824 10380 12880
rect 3988 12820 3994 12822
rect 5993 12819 6059 12822
rect 6310 12820 6316 12822
rect 6380 12822 10380 12824
rect 10504 12880 13511 12882
rect 10504 12824 13450 12880
rect 13506 12824 13511 12880
rect 10504 12822 13511 12824
rect 6380 12820 6427 12822
rect 6361 12819 6427 12820
rect 4337 12746 4403 12749
rect 4981 12746 5047 12749
rect 10504 12746 10564 12822
rect 13445 12819 13511 12822
rect 17493 12882 17559 12885
rect 19200 12882 20000 12912
rect 17493 12880 20000 12882
rect 17493 12824 17498 12880
rect 17554 12824 20000 12880
rect 17493 12822 20000 12824
rect 17493 12819 17559 12822
rect 19200 12792 20000 12822
rect 4337 12744 10564 12746
rect 4337 12688 4342 12744
rect 4398 12688 4986 12744
rect 5042 12688 10564 12744
rect 4337 12686 10564 12688
rect 11789 12746 11855 12749
rect 17585 12746 17651 12749
rect 11789 12744 17651 12746
rect 11789 12688 11794 12744
rect 11850 12688 17590 12744
rect 17646 12688 17651 12744
rect 11789 12686 17651 12688
rect 4337 12683 4403 12686
rect 4981 12683 5047 12686
rect 11789 12683 11855 12686
rect 17585 12683 17651 12686
rect 0 12610 800 12640
rect 2221 12610 2287 12613
rect 0 12608 2287 12610
rect 0 12552 2226 12608
rect 2282 12552 2287 12608
rect 0 12550 2287 12552
rect 0 12520 800 12550
rect 2221 12547 2287 12550
rect 3170 12544 3486 12545
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 16514 12479 16830 12480
rect 1710 12412 1716 12476
rect 1780 12474 1786 12476
rect 2957 12474 3023 12477
rect 1780 12472 3023 12474
rect 1780 12416 2962 12472
rect 3018 12416 3023 12472
rect 1780 12414 3023 12416
rect 1780 12412 1786 12414
rect 2957 12411 3023 12414
rect 12525 12474 12591 12477
rect 14549 12474 14615 12477
rect 12525 12472 14615 12474
rect 12525 12416 12530 12472
rect 12586 12416 14554 12472
rect 14610 12416 14615 12472
rect 12525 12414 14615 12416
rect 12525 12411 12591 12414
rect 14549 12411 14615 12414
rect 14958 12412 14964 12476
rect 15028 12474 15034 12476
rect 15101 12474 15167 12477
rect 15028 12472 15167 12474
rect 15028 12416 15106 12472
rect 15162 12416 15167 12472
rect 15028 12414 15167 12416
rect 15028 12412 15034 12414
rect 15101 12411 15167 12414
rect 17677 12474 17743 12477
rect 19200 12474 20000 12504
rect 17677 12472 20000 12474
rect 17677 12416 17682 12472
rect 17738 12416 20000 12472
rect 17677 12414 20000 12416
rect 17677 12411 17743 12414
rect 19200 12384 20000 12414
rect 1945 12338 2011 12341
rect 9673 12338 9739 12341
rect 13854 12338 13860 12340
rect 1945 12336 13860 12338
rect 1945 12280 1950 12336
rect 2006 12280 9678 12336
rect 9734 12280 13860 12336
rect 1945 12278 13860 12280
rect 1945 12275 2011 12278
rect 9673 12275 9739 12278
rect 13854 12276 13860 12278
rect 13924 12338 13930 12340
rect 15009 12338 15075 12341
rect 13924 12336 15075 12338
rect 13924 12280 15014 12336
rect 15070 12280 15075 12336
rect 13924 12278 15075 12280
rect 13924 12276 13930 12278
rect 15009 12275 15075 12278
rect 0 12202 800 12232
rect 2221 12202 2287 12205
rect 0 12200 2287 12202
rect 0 12144 2226 12200
rect 2282 12144 2287 12200
rect 0 12142 2287 12144
rect 0 12112 800 12142
rect 2221 12139 2287 12142
rect 3509 12202 3575 12205
rect 6545 12202 6611 12205
rect 13813 12202 13879 12205
rect 17953 12202 18019 12205
rect 3509 12200 6378 12202
rect 3509 12144 3514 12200
rect 3570 12144 6378 12200
rect 3509 12142 6378 12144
rect 3509 12139 3575 12142
rect 6318 12066 6378 12142
rect 6545 12200 13879 12202
rect 6545 12144 6550 12200
rect 6606 12144 13818 12200
rect 13874 12144 13879 12200
rect 6545 12142 13879 12144
rect 6545 12139 6611 12142
rect 13813 12139 13879 12142
rect 14046 12200 18019 12202
rect 14046 12144 17958 12200
rect 18014 12144 18019 12200
rect 14046 12142 18019 12144
rect 9397 12066 9463 12069
rect 6318 12064 9463 12066
rect 6318 12008 9402 12064
rect 9458 12008 9463 12064
rect 6318 12006 9463 12008
rect 9397 12003 9463 12006
rect 10409 12066 10475 12069
rect 14046 12066 14106 12142
rect 17953 12139 18019 12142
rect 10409 12064 14106 12066
rect 10409 12008 10414 12064
rect 10470 12008 14106 12064
rect 10409 12006 14106 12008
rect 16205 12066 16271 12069
rect 17677 12066 17743 12069
rect 19200 12066 20000 12096
rect 16205 12064 20000 12066
rect 16205 12008 16210 12064
rect 16266 12008 17682 12064
rect 17738 12008 20000 12064
rect 16205 12006 20000 12008
rect 10409 12003 10475 12006
rect 16205 12003 16271 12006
rect 17677 12003 17743 12006
rect 5394 12000 5710 12001
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 19200 11976 20000 12006
rect 14290 11935 14606 11936
rect 13486 11868 13492 11932
rect 13556 11930 13562 11932
rect 13813 11930 13879 11933
rect 13556 11928 13879 11930
rect 13556 11872 13818 11928
rect 13874 11872 13879 11928
rect 13556 11870 13879 11872
rect 13556 11868 13562 11870
rect 13813 11867 13879 11870
rect 0 11794 800 11824
rect 2037 11794 2103 11797
rect 0 11792 2103 11794
rect 0 11736 2042 11792
rect 2098 11736 2103 11792
rect 0 11734 2103 11736
rect 0 11704 800 11734
rect 2037 11731 2103 11734
rect 2773 11794 2839 11797
rect 3049 11794 3115 11797
rect 11789 11794 11855 11797
rect 2773 11792 11855 11794
rect 2773 11736 2778 11792
rect 2834 11736 3054 11792
rect 3110 11736 11794 11792
rect 11850 11736 11855 11792
rect 2773 11734 11855 11736
rect 2773 11731 2839 11734
rect 3049 11731 3115 11734
rect 11789 11731 11855 11734
rect 4981 11658 5047 11661
rect 9213 11658 9279 11661
rect 4981 11656 9279 11658
rect 4981 11600 4986 11656
rect 5042 11600 9218 11656
rect 9274 11600 9279 11656
rect 4981 11598 9279 11600
rect 4981 11595 5047 11598
rect 9213 11595 9279 11598
rect 9397 11658 9463 11661
rect 10777 11658 10843 11661
rect 9397 11656 10843 11658
rect 9397 11600 9402 11656
rect 9458 11600 10782 11656
rect 10838 11600 10843 11656
rect 9397 11598 10843 11600
rect 9397 11595 9463 11598
rect 10777 11595 10843 11598
rect 16389 11658 16455 11661
rect 18045 11658 18111 11661
rect 19200 11658 20000 11688
rect 16389 11656 20000 11658
rect 16389 11600 16394 11656
rect 16450 11600 18050 11656
rect 18106 11600 20000 11656
rect 16389 11598 20000 11600
rect 16389 11595 16455 11598
rect 18045 11595 18111 11598
rect 19200 11568 20000 11598
rect 9070 11460 9076 11524
rect 9140 11522 9146 11524
rect 9305 11522 9371 11525
rect 9140 11520 9371 11522
rect 9140 11464 9310 11520
rect 9366 11464 9371 11520
rect 9140 11462 9371 11464
rect 9140 11460 9146 11462
rect 9305 11459 9371 11462
rect 3170 11456 3486 11457
rect 0 11386 800 11416
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 16514 11391 16830 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 3785 11386 3851 11389
rect 4153 11386 4219 11389
rect 3785 11384 4219 11386
rect 3785 11328 3790 11384
rect 3846 11328 4158 11384
rect 4214 11328 4219 11384
rect 3785 11326 4219 11328
rect 3785 11323 3851 11326
rect 4153 11323 4219 11326
rect 5022 11324 5028 11388
rect 5092 11386 5098 11388
rect 5809 11386 5875 11389
rect 5092 11384 5875 11386
rect 5092 11328 5814 11384
rect 5870 11328 5875 11384
rect 5092 11326 5875 11328
rect 5092 11324 5098 11326
rect 5809 11323 5875 11326
rect 2497 11250 2563 11253
rect 10225 11250 10291 11253
rect 2497 11248 10291 11250
rect 2497 11192 2502 11248
rect 2558 11192 10230 11248
rect 10286 11192 10291 11248
rect 2497 11190 10291 11192
rect 2497 11187 2563 11190
rect 10225 11187 10291 11190
rect 10409 11250 10475 11253
rect 14549 11250 14615 11253
rect 10409 11248 14615 11250
rect 10409 11192 10414 11248
rect 10470 11192 14554 11248
rect 14610 11192 14615 11248
rect 10409 11190 14615 11192
rect 10409 11187 10475 11190
rect 14549 11187 14615 11190
rect 18413 11250 18479 11253
rect 19200 11250 20000 11280
rect 18413 11248 20000 11250
rect 18413 11192 18418 11248
rect 18474 11192 20000 11248
rect 18413 11190 20000 11192
rect 18413 11187 18479 11190
rect 19200 11160 20000 11190
rect 1945 11114 2011 11117
rect 4981 11114 5047 11117
rect 1945 11112 5047 11114
rect 1945 11056 1950 11112
rect 2006 11056 4986 11112
rect 5042 11056 5047 11112
rect 1945 11054 5047 11056
rect 1945 11051 2011 11054
rect 4981 11051 5047 11054
rect 5206 11052 5212 11116
rect 5276 11114 5282 11116
rect 6821 11114 6887 11117
rect 5276 11112 6887 11114
rect 5276 11056 6826 11112
rect 6882 11056 6887 11112
rect 5276 11054 6887 11056
rect 5276 11052 5282 11054
rect 6821 11051 6887 11054
rect 7189 11114 7255 11117
rect 9213 11116 9279 11117
rect 7414 11114 7420 11116
rect 7189 11112 7420 11114
rect 7189 11056 7194 11112
rect 7250 11056 7420 11112
rect 7189 11054 7420 11056
rect 7189 11051 7255 11054
rect 7414 11052 7420 11054
rect 7484 11052 7490 11116
rect 9213 11114 9260 11116
rect 9168 11112 9260 11114
rect 9168 11056 9218 11112
rect 9168 11054 9260 11056
rect 9213 11052 9260 11054
rect 9324 11052 9330 11116
rect 14089 11114 14155 11117
rect 15745 11114 15811 11117
rect 14089 11112 15811 11114
rect 14089 11056 14094 11112
rect 14150 11056 15750 11112
rect 15806 11056 15811 11112
rect 14089 11054 15811 11056
rect 9213 11051 9279 11052
rect 14089 11051 14155 11054
rect 15745 11051 15811 11054
rect 16757 11114 16823 11117
rect 17585 11114 17651 11117
rect 17861 11114 17927 11117
rect 16757 11112 17927 11114
rect 16757 11056 16762 11112
rect 16818 11056 17590 11112
rect 17646 11056 17866 11112
rect 17922 11056 17927 11112
rect 16757 11054 17927 11056
rect 16757 11051 16823 11054
rect 17585 11051 17651 11054
rect 17861 11051 17927 11054
rect 0 10978 800 11008
rect 2221 10978 2287 10981
rect 0 10976 2287 10978
rect 0 10920 2226 10976
rect 2282 10920 2287 10976
rect 0 10918 2287 10920
rect 0 10888 800 10918
rect 2221 10915 2287 10918
rect 2405 10978 2471 10981
rect 4981 10978 5047 10981
rect 2405 10976 5047 10978
rect 2405 10920 2410 10976
rect 2466 10920 4986 10976
rect 5042 10920 5047 10976
rect 2405 10918 5047 10920
rect 2405 10915 2471 10918
rect 4981 10915 5047 10918
rect 15929 10978 15995 10981
rect 16849 10978 16915 10981
rect 15929 10976 16915 10978
rect 15929 10920 15934 10976
rect 15990 10920 16854 10976
rect 16910 10920 16915 10976
rect 15929 10918 16915 10920
rect 15929 10915 15995 10918
rect 16849 10915 16915 10918
rect 17033 10978 17099 10981
rect 18505 10978 18571 10981
rect 17033 10976 18571 10978
rect 17033 10920 17038 10976
rect 17094 10920 18510 10976
rect 18566 10920 18571 10976
rect 17033 10918 18571 10920
rect 17033 10915 17099 10918
rect 18505 10915 18571 10918
rect 5394 10912 5710 10913
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 14290 10847 14606 10848
rect 3969 10844 4035 10845
rect 3918 10780 3924 10844
rect 3988 10842 4035 10844
rect 4981 10842 5047 10845
rect 3988 10840 5047 10842
rect 4030 10784 4986 10840
rect 5042 10784 5047 10840
rect 3988 10782 5047 10784
rect 3988 10780 4035 10782
rect 3969 10779 4035 10780
rect 4981 10779 5047 10782
rect 5809 10842 5875 10845
rect 9029 10842 9095 10845
rect 5809 10840 9095 10842
rect 5809 10784 5814 10840
rect 5870 10784 9034 10840
rect 9090 10784 9095 10840
rect 5809 10782 9095 10784
rect 5809 10779 5875 10782
rect 9029 10779 9095 10782
rect 14733 10842 14799 10845
rect 16941 10842 17007 10845
rect 14733 10840 17007 10842
rect 14733 10784 14738 10840
rect 14794 10784 16946 10840
rect 17002 10784 17007 10840
rect 14733 10782 17007 10784
rect 14733 10779 14799 10782
rect 16941 10779 17007 10782
rect 17677 10842 17743 10845
rect 19200 10842 20000 10872
rect 17677 10840 20000 10842
rect 17677 10784 17682 10840
rect 17738 10784 20000 10840
rect 17677 10782 20000 10784
rect 17677 10779 17743 10782
rect 19200 10752 20000 10782
rect 2814 10644 2820 10708
rect 2884 10706 2890 10708
rect 3049 10706 3115 10709
rect 2884 10704 3115 10706
rect 2884 10648 3054 10704
rect 3110 10648 3115 10704
rect 2884 10646 3115 10648
rect 2884 10644 2890 10646
rect 3049 10643 3115 10646
rect 3601 10706 3667 10709
rect 11329 10706 11395 10709
rect 3601 10704 11395 10706
rect 3601 10648 3606 10704
rect 3662 10648 11334 10704
rect 11390 10648 11395 10704
rect 3601 10646 11395 10648
rect 3601 10643 3667 10646
rect 11329 10643 11395 10646
rect 11697 10706 11763 10709
rect 17953 10706 18019 10709
rect 11697 10704 18019 10706
rect 11697 10648 11702 10704
rect 11758 10648 17958 10704
rect 18014 10648 18019 10704
rect 11697 10646 18019 10648
rect 11697 10643 11763 10646
rect 17953 10643 18019 10646
rect 0 10570 800 10600
rect 1485 10570 1551 10573
rect 0 10568 1551 10570
rect 0 10512 1490 10568
rect 1546 10512 1551 10568
rect 0 10510 1551 10512
rect 0 10480 800 10510
rect 1485 10507 1551 10510
rect 4981 10570 5047 10573
rect 18045 10570 18111 10573
rect 4981 10568 18111 10570
rect 4981 10512 4986 10568
rect 5042 10512 18050 10568
rect 18106 10512 18111 10568
rect 4981 10510 18111 10512
rect 4981 10507 5047 10510
rect 18045 10507 18111 10510
rect 3601 10434 3667 10437
rect 4613 10434 4679 10437
rect 5165 10434 5231 10437
rect 3601 10432 4679 10434
rect 3601 10376 3606 10432
rect 3662 10376 4618 10432
rect 4674 10376 4679 10432
rect 3601 10374 4679 10376
rect 3601 10371 3667 10374
rect 4613 10371 4679 10374
rect 4984 10432 5231 10434
rect 4984 10376 5170 10432
rect 5226 10376 5231 10432
rect 4984 10374 5231 10376
rect 3170 10368 3486 10369
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 4984 10301 5044 10374
rect 5165 10371 5231 10374
rect 6361 10434 6427 10437
rect 6494 10434 6500 10436
rect 6361 10432 6500 10434
rect 6361 10376 6366 10432
rect 6422 10376 6500 10432
rect 6361 10374 6500 10376
rect 6361 10371 6427 10374
rect 6494 10372 6500 10374
rect 6564 10372 6570 10436
rect 16982 10372 16988 10436
rect 17052 10434 17058 10436
rect 17861 10434 17927 10437
rect 17052 10432 17927 10434
rect 17052 10376 17866 10432
rect 17922 10376 17927 10432
rect 17052 10374 17927 10376
rect 17052 10372 17058 10374
rect 17861 10371 17927 10374
rect 18413 10434 18479 10437
rect 19200 10434 20000 10464
rect 18413 10432 20000 10434
rect 18413 10376 18418 10432
rect 18474 10376 20000 10432
rect 18413 10374 20000 10376
rect 18413 10371 18479 10374
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 19200 10344 20000 10374
rect 16514 10303 16830 10304
rect 4981 10296 5047 10301
rect 4981 10240 4986 10296
rect 5042 10240 5047 10296
rect 4981 10235 5047 10240
rect 5257 10298 5323 10301
rect 5942 10298 5948 10300
rect 5257 10296 5948 10298
rect 5257 10240 5262 10296
rect 5318 10240 5948 10296
rect 5257 10238 5948 10240
rect 5257 10235 5323 10238
rect 5942 10236 5948 10238
rect 6012 10236 6018 10300
rect 15561 10298 15627 10301
rect 16062 10298 16068 10300
rect 15561 10296 16068 10298
rect 15561 10240 15566 10296
rect 15622 10240 16068 10296
rect 15561 10238 16068 10240
rect 15561 10235 15627 10238
rect 16062 10236 16068 10238
rect 16132 10236 16138 10300
rect 0 10162 800 10192
rect 3049 10162 3115 10165
rect 11421 10162 11487 10165
rect 12433 10162 12499 10165
rect 18321 10162 18387 10165
rect 0 10102 1410 10162
rect 0 10072 800 10102
rect 1350 9890 1410 10102
rect 3049 10160 18387 10162
rect 3049 10104 3054 10160
rect 3110 10104 11426 10160
rect 11482 10104 12438 10160
rect 12494 10104 18326 10160
rect 18382 10104 18387 10160
rect 3049 10102 18387 10104
rect 3049 10099 3115 10102
rect 11421 10099 11487 10102
rect 12433 10099 12499 10102
rect 18321 10099 18387 10102
rect 1669 10026 1735 10029
rect 4245 10026 4311 10029
rect 1669 10024 4311 10026
rect 1669 9968 1674 10024
rect 1730 9968 4250 10024
rect 4306 9968 4311 10024
rect 1669 9966 4311 9968
rect 1669 9963 1735 9966
rect 4245 9963 4311 9966
rect 4470 9964 4476 10028
rect 4540 10026 4546 10028
rect 5441 10026 5507 10029
rect 4540 10024 5507 10026
rect 4540 9968 5446 10024
rect 5502 9968 5507 10024
rect 4540 9966 5507 9968
rect 4540 9964 4546 9966
rect 5441 9963 5507 9966
rect 5717 10026 5783 10029
rect 11697 10026 11763 10029
rect 5717 10024 11763 10026
rect 5717 9968 5722 10024
rect 5778 9968 11702 10024
rect 11758 9968 11763 10024
rect 5717 9966 11763 9968
rect 5717 9963 5783 9966
rect 11697 9963 11763 9966
rect 11881 10026 11947 10029
rect 15929 10026 15995 10029
rect 16113 10028 16179 10029
rect 11881 10024 15995 10026
rect 11881 9968 11886 10024
rect 11942 9968 15934 10024
rect 15990 9968 15995 10024
rect 11881 9966 15995 9968
rect 11881 9963 11947 9966
rect 15929 9963 15995 9966
rect 16062 9964 16068 10028
rect 16132 10026 16179 10028
rect 16389 10026 16455 10029
rect 19200 10026 20000 10056
rect 16132 10024 16224 10026
rect 16174 9968 16224 10024
rect 16132 9966 16224 9968
rect 16389 10024 20000 10026
rect 16389 9968 16394 10024
rect 16450 9968 20000 10024
rect 16389 9966 20000 9968
rect 16132 9964 16179 9966
rect 16113 9963 16179 9964
rect 16389 9963 16455 9966
rect 19200 9936 20000 9966
rect 1485 9890 1551 9893
rect 1350 9888 1551 9890
rect 1350 9832 1490 9888
rect 1546 9832 1551 9888
rect 1350 9830 1551 9832
rect 1485 9827 1551 9830
rect 3509 9890 3575 9893
rect 4889 9890 4955 9893
rect 3509 9888 4955 9890
rect 3509 9832 3514 9888
rect 3570 9832 4894 9888
rect 4950 9832 4955 9888
rect 3509 9830 4955 9832
rect 3509 9827 3575 9830
rect 4889 9827 4955 9830
rect 6821 9890 6887 9893
rect 7465 9890 7531 9893
rect 6821 9888 7531 9890
rect 6821 9832 6826 9888
rect 6882 9832 7470 9888
rect 7526 9832 7531 9888
rect 6821 9830 7531 9832
rect 6821 9827 6887 9830
rect 7465 9827 7531 9830
rect 15285 9890 15351 9893
rect 16481 9890 16547 9893
rect 17033 9892 17099 9893
rect 15285 9888 16547 9890
rect 15285 9832 15290 9888
rect 15346 9832 16486 9888
rect 16542 9832 16547 9888
rect 15285 9830 16547 9832
rect 15285 9827 15351 9830
rect 16481 9827 16547 9830
rect 16982 9828 16988 9892
rect 17052 9890 17099 9892
rect 17052 9888 17144 9890
rect 17094 9832 17144 9888
rect 17052 9830 17144 9832
rect 17052 9828 17099 9830
rect 17033 9827 17099 9828
rect 5394 9824 5710 9825
rect 0 9754 800 9784
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 14290 9759 14606 9760
rect 2221 9754 2287 9757
rect 0 9752 2287 9754
rect 0 9696 2226 9752
rect 2282 9696 2287 9752
rect 0 9694 2287 9696
rect 0 9664 800 9694
rect 2221 9691 2287 9694
rect 2865 9754 2931 9757
rect 2998 9754 3004 9756
rect 2865 9752 3004 9754
rect 2865 9696 2870 9752
rect 2926 9696 3004 9752
rect 2865 9694 3004 9696
rect 2865 9691 2931 9694
rect 2998 9692 3004 9694
rect 3068 9692 3074 9756
rect 3969 9754 4035 9757
rect 4102 9754 4108 9756
rect 3969 9752 4108 9754
rect 3969 9696 3974 9752
rect 4030 9696 4108 9752
rect 3969 9694 4108 9696
rect 3969 9691 4035 9694
rect 4102 9692 4108 9694
rect 4172 9692 4178 9756
rect 6637 9754 6703 9757
rect 6862 9754 6868 9756
rect 6637 9752 6868 9754
rect 6637 9696 6642 9752
rect 6698 9696 6868 9752
rect 6637 9694 6868 9696
rect 6637 9691 6703 9694
rect 6862 9692 6868 9694
rect 6932 9692 6938 9756
rect 7925 9754 7991 9757
rect 13997 9756 14063 9757
rect 8150 9754 8156 9756
rect 7925 9752 8156 9754
rect 7925 9696 7930 9752
rect 7986 9696 8156 9752
rect 7925 9694 8156 9696
rect 7925 9691 7991 9694
rect 8150 9692 8156 9694
rect 8220 9692 8226 9756
rect 13997 9752 14044 9756
rect 14108 9754 14114 9756
rect 14733 9754 14799 9757
rect 16941 9754 17007 9757
rect 13997 9696 14002 9752
rect 13997 9692 14044 9696
rect 14108 9694 14154 9754
rect 14733 9752 17007 9754
rect 14733 9696 14738 9752
rect 14794 9696 16946 9752
rect 17002 9696 17007 9752
rect 14733 9694 17007 9696
rect 14108 9692 14114 9694
rect 13997 9691 14063 9692
rect 14733 9691 14799 9694
rect 16941 9691 17007 9694
rect 17861 9756 17927 9757
rect 17861 9752 17908 9756
rect 17972 9754 17978 9756
rect 17861 9696 17866 9752
rect 17861 9692 17908 9696
rect 17972 9694 18018 9754
rect 17972 9692 17978 9694
rect 17861 9691 17927 9692
rect 3049 9618 3115 9621
rect 7833 9618 7899 9621
rect 3049 9616 3986 9618
rect 3049 9560 3054 9616
rect 3110 9560 3986 9616
rect 3049 9558 3986 9560
rect 3049 9555 3115 9558
rect 3601 9482 3667 9485
rect 3734 9482 3740 9484
rect 3601 9480 3740 9482
rect 3601 9424 3606 9480
rect 3662 9424 3740 9480
rect 3601 9422 3740 9424
rect 3601 9419 3667 9422
rect 3734 9420 3740 9422
rect 3804 9420 3810 9484
rect 0 9346 800 9376
rect 2865 9346 2931 9349
rect 0 9344 2931 9346
rect 0 9288 2870 9344
rect 2926 9288 2931 9344
rect 0 9286 2931 9288
rect 0 9256 800 9286
rect 2865 9283 2931 9286
rect 3170 9280 3486 9281
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 3926 9210 3986 9558
rect 5030 9616 7899 9618
rect 5030 9560 7838 9616
rect 7894 9560 7899 9616
rect 5030 9558 7899 9560
rect 4521 9482 4587 9485
rect 4654 9482 4660 9484
rect 4521 9480 4660 9482
rect 4521 9424 4526 9480
rect 4582 9424 4660 9480
rect 4521 9422 4660 9424
rect 4521 9419 4587 9422
rect 4654 9420 4660 9422
rect 4724 9420 4730 9484
rect 4153 9346 4219 9349
rect 5030 9346 5090 9558
rect 7833 9555 7899 9558
rect 8661 9618 8727 9621
rect 16021 9618 16087 9621
rect 8661 9616 16087 9618
rect 8661 9560 8666 9616
rect 8722 9560 16026 9616
rect 16082 9560 16087 9616
rect 8661 9558 16087 9560
rect 8661 9555 8727 9558
rect 13310 9485 13370 9558
rect 16021 9555 16087 9558
rect 16297 9618 16363 9621
rect 19200 9618 20000 9648
rect 16297 9616 20000 9618
rect 16297 9560 16302 9616
rect 16358 9560 20000 9616
rect 16297 9558 20000 9560
rect 16297 9555 16363 9558
rect 19200 9528 20000 9558
rect 5942 9420 5948 9484
rect 6012 9482 6018 9484
rect 10225 9482 10291 9485
rect 6012 9480 10291 9482
rect 6012 9424 10230 9480
rect 10286 9424 10291 9480
rect 6012 9422 10291 9424
rect 6012 9420 6018 9422
rect 10225 9419 10291 9422
rect 13261 9480 13370 9485
rect 13261 9424 13266 9480
rect 13322 9424 13370 9480
rect 13261 9422 13370 9424
rect 16205 9482 16271 9485
rect 16205 9480 17050 9482
rect 16205 9424 16210 9480
rect 16266 9424 17050 9480
rect 16205 9422 17050 9424
rect 13261 9419 13327 9422
rect 16205 9419 16271 9422
rect 4153 9344 5090 9346
rect 4153 9288 4158 9344
rect 4214 9288 5090 9344
rect 4153 9286 5090 9288
rect 5993 9346 6059 9349
rect 6361 9346 6427 9349
rect 5993 9344 6427 9346
rect 5993 9288 5998 9344
rect 6054 9288 6366 9344
rect 6422 9288 6427 9344
rect 5993 9286 6427 9288
rect 4153 9283 4219 9286
rect 5993 9283 6059 9286
rect 6361 9283 6427 9286
rect 13486 9284 13492 9348
rect 13556 9346 13562 9348
rect 14365 9346 14431 9349
rect 14825 9348 14891 9349
rect 13556 9344 14431 9346
rect 13556 9288 14370 9344
rect 14426 9288 14431 9344
rect 13556 9286 14431 9288
rect 13556 9284 13562 9286
rect 14365 9283 14431 9286
rect 14774 9284 14780 9348
rect 14844 9346 14891 9348
rect 14844 9344 14936 9346
rect 14886 9288 14936 9344
rect 14844 9286 14936 9288
rect 14844 9284 14891 9286
rect 14825 9283 14891 9284
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 16514 9215 16830 9216
rect 5901 9210 5967 9213
rect 13445 9210 13511 9213
rect 14181 9210 14247 9213
rect 3926 9208 7482 9210
rect 3926 9152 5906 9208
rect 5962 9152 7482 9208
rect 3926 9150 7482 9152
rect 5901 9147 5967 9150
rect 3325 9074 3391 9077
rect 4470 9074 4476 9076
rect 3325 9072 4476 9074
rect 3325 9016 3330 9072
rect 3386 9016 4476 9072
rect 3325 9014 4476 9016
rect 3325 9011 3391 9014
rect 4470 9012 4476 9014
rect 4540 9012 4546 9076
rect 5625 9074 5691 9077
rect 6269 9074 6335 9077
rect 5625 9072 6335 9074
rect 5625 9016 5630 9072
rect 5686 9016 6274 9072
rect 6330 9016 6335 9072
rect 5625 9014 6335 9016
rect 7422 9074 7482 9150
rect 13445 9208 14247 9210
rect 13445 9152 13450 9208
rect 13506 9152 14186 9208
rect 14242 9152 14247 9208
rect 13445 9150 14247 9152
rect 13445 9147 13511 9150
rect 14181 9147 14247 9150
rect 14457 9210 14523 9213
rect 15745 9210 15811 9213
rect 14457 9208 15811 9210
rect 14457 9152 14462 9208
rect 14518 9152 15750 9208
rect 15806 9152 15811 9208
rect 14457 9150 15811 9152
rect 14457 9147 14523 9150
rect 15745 9147 15811 9150
rect 15929 9210 15995 9213
rect 16297 9210 16363 9213
rect 15929 9208 16363 9210
rect 15929 9152 15934 9208
rect 15990 9152 16302 9208
rect 16358 9152 16363 9208
rect 15929 9150 16363 9152
rect 16990 9210 17050 9422
rect 19200 9210 20000 9240
rect 16990 9150 20000 9210
rect 15929 9147 15995 9150
rect 16297 9147 16363 9150
rect 19200 9120 20000 9150
rect 8569 9074 8635 9077
rect 7422 9072 8635 9074
rect 7422 9016 8574 9072
rect 8630 9016 8635 9072
rect 7422 9014 8635 9016
rect 5625 9011 5691 9014
rect 6269 9011 6335 9014
rect 8569 9011 8635 9014
rect 9765 9074 9831 9077
rect 11329 9074 11395 9077
rect 9765 9072 11395 9074
rect 9765 9016 9770 9072
rect 9826 9016 11334 9072
rect 11390 9016 11395 9072
rect 9765 9014 11395 9016
rect 9765 9011 9831 9014
rect 11329 9011 11395 9014
rect 11789 9074 11855 9077
rect 14825 9074 14891 9077
rect 17677 9074 17743 9077
rect 11789 9072 17743 9074
rect 11789 9016 11794 9072
rect 11850 9016 14830 9072
rect 14886 9016 17682 9072
rect 17738 9016 17743 9072
rect 11789 9014 17743 9016
rect 11789 9011 11855 9014
rect 14825 9011 14891 9014
rect 17677 9011 17743 9014
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 2405 8940 2471 8941
rect 2405 8938 2452 8940
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 2360 8936 2452 8938
rect 2360 8880 2410 8936
rect 2360 8878 2452 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 2405 8876 2452 8878
rect 2516 8876 2522 8940
rect 5809 8938 5875 8941
rect 16205 8938 16271 8941
rect 5809 8936 16271 8938
rect 5809 8880 5814 8936
rect 5870 8880 16210 8936
rect 16266 8880 16271 8936
rect 5809 8878 16271 8880
rect 2405 8875 2471 8876
rect 5809 8875 5875 8878
rect 16205 8875 16271 8878
rect 1761 8802 1827 8805
rect 1894 8802 1900 8804
rect 1761 8800 1900 8802
rect 1761 8744 1766 8800
rect 1822 8744 1900 8800
rect 1761 8742 1900 8744
rect 1761 8739 1827 8742
rect 1894 8740 1900 8742
rect 1964 8740 1970 8804
rect 3785 8802 3851 8805
rect 5022 8802 5028 8804
rect 2086 8800 5028 8802
rect 2086 8744 3790 8800
rect 3846 8744 5028 8800
rect 2086 8742 5028 8744
rect 1761 8666 1827 8669
rect 2086 8666 2146 8742
rect 3785 8739 3851 8742
rect 5022 8740 5028 8742
rect 5092 8740 5098 8804
rect 15193 8802 15259 8805
rect 19200 8802 20000 8832
rect 15193 8800 20000 8802
rect 15193 8744 15198 8800
rect 15254 8744 20000 8800
rect 15193 8742 20000 8744
rect 15193 8739 15259 8742
rect 5394 8736 5710 8737
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 19200 8712 20000 8742
rect 14290 8671 14606 8672
rect 1761 8664 2146 8666
rect 1761 8608 1766 8664
rect 1822 8608 2146 8664
rect 1761 8606 2146 8608
rect 2313 8666 2379 8669
rect 4153 8666 4219 8669
rect 2313 8664 4219 8666
rect 2313 8608 2318 8664
rect 2374 8608 4158 8664
rect 4214 8608 4219 8664
rect 2313 8606 4219 8608
rect 1761 8603 1827 8606
rect 2313 8603 2379 8606
rect 4153 8603 4219 8606
rect 13629 8666 13695 8669
rect 13854 8666 13860 8668
rect 13629 8664 13860 8666
rect 13629 8608 13634 8664
rect 13690 8608 13860 8664
rect 13629 8606 13860 8608
rect 13629 8603 13695 8606
rect 13854 8604 13860 8606
rect 13924 8604 13930 8668
rect 14733 8666 14799 8669
rect 18045 8666 18111 8669
rect 14733 8664 18111 8666
rect 14733 8608 14738 8664
rect 14794 8608 18050 8664
rect 18106 8608 18111 8664
rect 14733 8606 18111 8608
rect 14733 8603 14799 8606
rect 18045 8603 18111 8606
rect 0 8530 800 8560
rect 2957 8530 3023 8533
rect 0 8528 3023 8530
rect 0 8472 2962 8528
rect 3018 8472 3023 8528
rect 0 8470 3023 8472
rect 0 8440 800 8470
rect 2957 8467 3023 8470
rect 3877 8530 3943 8533
rect 9489 8530 9555 8533
rect 3877 8528 9555 8530
rect 3877 8472 3882 8528
rect 3938 8472 9494 8528
rect 9550 8472 9555 8528
rect 3877 8470 9555 8472
rect 3877 8467 3943 8470
rect 9489 8467 9555 8470
rect 13353 8530 13419 8533
rect 13353 8528 15762 8530
rect 13353 8472 13358 8528
rect 13414 8472 15762 8528
rect 13353 8470 15762 8472
rect 13353 8467 13419 8470
rect 1301 8394 1367 8397
rect 3417 8394 3483 8397
rect 1301 8392 3483 8394
rect 1301 8336 1306 8392
rect 1362 8336 3422 8392
rect 3478 8336 3483 8392
rect 1301 8334 3483 8336
rect 1301 8331 1367 8334
rect 3417 8331 3483 8334
rect 8017 8394 8083 8397
rect 11605 8394 11671 8397
rect 15561 8394 15627 8397
rect 8017 8392 15627 8394
rect 8017 8336 8022 8392
rect 8078 8336 11610 8392
rect 11666 8336 15566 8392
rect 15622 8336 15627 8392
rect 8017 8334 15627 8336
rect 15702 8394 15762 8470
rect 16757 8394 16823 8397
rect 17493 8394 17559 8397
rect 15702 8392 17559 8394
rect 15702 8336 16762 8392
rect 16818 8336 17498 8392
rect 17554 8336 17559 8392
rect 15702 8334 17559 8336
rect 8017 8331 8083 8334
rect 11605 8331 11671 8334
rect 15561 8331 15627 8334
rect 16757 8331 16823 8334
rect 17493 8331 17559 8334
rect 18413 8394 18479 8397
rect 19200 8394 20000 8424
rect 18413 8392 20000 8394
rect 18413 8336 18418 8392
rect 18474 8336 20000 8392
rect 18413 8334 20000 8336
rect 18413 8331 18479 8334
rect 19200 8304 20000 8334
rect 6545 8260 6611 8261
rect 6494 8258 6500 8260
rect 6454 8198 6500 8258
rect 6564 8256 6611 8260
rect 6606 8200 6611 8256
rect 6494 8196 6500 8198
rect 6564 8196 6611 8200
rect 6545 8195 6611 8196
rect 3170 8192 3486 8193
rect 0 8122 800 8152
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 16514 8127 16830 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 13997 8122 14063 8125
rect 13997 8120 16314 8122
rect 13997 8064 14002 8120
rect 14058 8064 16314 8120
rect 13997 8062 16314 8064
rect 13997 8059 14063 8062
rect 2037 7986 2103 7989
rect 3601 7986 3667 7989
rect 2037 7984 3667 7986
rect 2037 7928 2042 7984
rect 2098 7928 3606 7984
rect 3662 7928 3667 7984
rect 2037 7926 3667 7928
rect 2037 7923 2103 7926
rect 3601 7923 3667 7926
rect 4153 7986 4219 7989
rect 9305 7986 9371 7989
rect 4153 7984 9371 7986
rect 4153 7928 4158 7984
rect 4214 7928 9310 7984
rect 9366 7928 9371 7984
rect 4153 7926 9371 7928
rect 4153 7923 4219 7926
rect 9305 7923 9371 7926
rect 10225 7986 10291 7989
rect 15193 7986 15259 7989
rect 10225 7984 15259 7986
rect 10225 7928 10230 7984
rect 10286 7928 15198 7984
rect 15254 7928 15259 7984
rect 10225 7926 15259 7928
rect 16254 7986 16314 8062
rect 16757 7986 16823 7989
rect 16254 7984 16823 7986
rect 16254 7928 16762 7984
rect 16818 7928 16823 7984
rect 16254 7926 16823 7928
rect 10225 7923 10291 7926
rect 15193 7923 15259 7926
rect 16757 7923 16823 7926
rect 18505 7986 18571 7989
rect 19200 7986 20000 8016
rect 18505 7984 20000 7986
rect 18505 7928 18510 7984
rect 18566 7928 20000 7984
rect 18505 7926 20000 7928
rect 18505 7923 18571 7926
rect 19200 7896 20000 7926
rect 5073 7850 5139 7853
rect 5717 7850 5783 7853
rect 12985 7850 13051 7853
rect 5073 7848 13051 7850
rect 5073 7792 5078 7848
rect 5134 7792 5722 7848
rect 5778 7792 12990 7848
rect 13046 7792 13051 7848
rect 5073 7790 13051 7792
rect 5073 7787 5139 7790
rect 5717 7787 5783 7790
rect 12985 7787 13051 7790
rect 13629 7850 13695 7853
rect 17953 7850 18019 7853
rect 13629 7848 18019 7850
rect 13629 7792 13634 7848
rect 13690 7792 17958 7848
rect 18014 7792 18019 7848
rect 13629 7790 18019 7792
rect 13629 7787 13695 7790
rect 17953 7787 18019 7790
rect 0 7714 800 7744
rect 1853 7714 1919 7717
rect 0 7712 1919 7714
rect 0 7656 1858 7712
rect 1914 7656 1919 7712
rect 0 7654 1919 7656
rect 0 7624 800 7654
rect 1853 7651 1919 7654
rect 14825 7714 14891 7717
rect 17493 7714 17559 7717
rect 14825 7712 17559 7714
rect 14825 7656 14830 7712
rect 14886 7656 17498 7712
rect 17554 7656 17559 7712
rect 14825 7654 17559 7656
rect 14825 7651 14891 7654
rect 17493 7651 17559 7654
rect 5394 7648 5710 7649
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 14290 7583 14606 7584
rect 4337 7578 4403 7581
rect 5206 7578 5212 7580
rect 2730 7576 5212 7578
rect 2730 7520 4342 7576
rect 4398 7520 5212 7576
rect 2730 7518 5212 7520
rect 2221 7442 2287 7445
rect 2730 7442 2790 7518
rect 4337 7515 4403 7518
rect 5206 7516 5212 7518
rect 5276 7516 5282 7580
rect 13629 7578 13695 7581
rect 12390 7576 13695 7578
rect 12390 7520 13634 7576
rect 13690 7520 13695 7576
rect 12390 7518 13695 7520
rect 2221 7440 2790 7442
rect 2221 7384 2226 7440
rect 2282 7384 2790 7440
rect 2221 7382 2790 7384
rect 2221 7379 2287 7382
rect 3734 7380 3740 7444
rect 3804 7442 3810 7444
rect 4061 7442 4127 7445
rect 3804 7440 4127 7442
rect 3804 7384 4066 7440
rect 4122 7384 4127 7440
rect 3804 7382 4127 7384
rect 3804 7380 3810 7382
rect 4061 7379 4127 7382
rect 4429 7442 4495 7445
rect 5533 7442 5599 7445
rect 6310 7442 6316 7444
rect 4429 7440 6316 7442
rect 4429 7384 4434 7440
rect 4490 7384 5538 7440
rect 5594 7384 6316 7440
rect 4429 7382 6316 7384
rect 4429 7379 4495 7382
rect 5533 7379 5599 7382
rect 6310 7380 6316 7382
rect 6380 7380 6386 7444
rect 9254 7380 9260 7444
rect 9324 7442 9330 7444
rect 12390 7442 12450 7518
rect 13629 7515 13695 7518
rect 18045 7578 18111 7581
rect 19200 7578 20000 7608
rect 18045 7576 20000 7578
rect 18045 7520 18050 7576
rect 18106 7520 20000 7576
rect 18045 7518 20000 7520
rect 18045 7515 18111 7518
rect 19200 7488 20000 7518
rect 9324 7382 12450 7442
rect 12893 7442 12959 7445
rect 16849 7442 16915 7445
rect 12893 7440 16915 7442
rect 12893 7384 12898 7440
rect 12954 7384 16854 7440
rect 16910 7384 16915 7440
rect 12893 7382 16915 7384
rect 9324 7380 9330 7382
rect 12893 7379 12959 7382
rect 16849 7379 16915 7382
rect 0 7306 800 7336
rect 1485 7306 1551 7309
rect 0 7304 1551 7306
rect 0 7248 1490 7304
rect 1546 7248 1551 7304
rect 0 7246 1551 7248
rect 0 7216 800 7246
rect 1485 7243 1551 7246
rect 2446 7244 2452 7308
rect 2516 7306 2522 7308
rect 3141 7306 3207 7309
rect 11697 7306 11763 7309
rect 2516 7304 11763 7306
rect 2516 7248 3146 7304
rect 3202 7248 11702 7304
rect 11758 7248 11763 7304
rect 2516 7246 11763 7248
rect 2516 7244 2522 7246
rect 3141 7243 3207 7246
rect 11697 7243 11763 7246
rect 13537 7306 13603 7309
rect 17125 7306 17191 7309
rect 13537 7304 17191 7306
rect 13537 7248 13542 7304
rect 13598 7248 17130 7304
rect 17186 7248 17191 7304
rect 13537 7246 17191 7248
rect 13537 7243 13603 7246
rect 17125 7243 17191 7246
rect 18413 7170 18479 7173
rect 19200 7170 20000 7200
rect 18413 7168 20000 7170
rect 18413 7112 18418 7168
rect 18474 7112 20000 7168
rect 18413 7110 20000 7112
rect 18413 7107 18479 7110
rect 3170 7104 3486 7105
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 19200 7080 20000 7110
rect 16514 7039 16830 7040
rect 17769 7036 17835 7037
rect 17718 7034 17724 7036
rect 17678 6974 17724 7034
rect 17788 7032 17835 7036
rect 17830 6976 17835 7032
rect 17718 6972 17724 6974
rect 17788 6972 17835 6976
rect 17769 6971 17835 6972
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 2497 6898 2563 6901
rect 5717 6898 5783 6901
rect 2497 6896 5783 6898
rect 2497 6840 2502 6896
rect 2558 6840 5722 6896
rect 5778 6840 5783 6896
rect 2497 6838 5783 6840
rect 2497 6835 2563 6838
rect 5717 6835 5783 6838
rect 12985 6898 13051 6901
rect 16665 6898 16731 6901
rect 12985 6896 16731 6898
rect 12985 6840 12990 6896
rect 13046 6840 16670 6896
rect 16726 6840 16731 6896
rect 12985 6838 16731 6840
rect 12985 6835 13051 6838
rect 16665 6835 16731 6838
rect 3325 6762 3391 6765
rect 3550 6762 3556 6764
rect 3325 6760 3556 6762
rect 3325 6704 3330 6760
rect 3386 6704 3556 6760
rect 3325 6702 3556 6704
rect 3325 6699 3391 6702
rect 3550 6700 3556 6702
rect 3620 6762 3626 6764
rect 4153 6762 4219 6765
rect 3620 6760 4219 6762
rect 3620 6704 4158 6760
rect 4214 6704 4219 6760
rect 3620 6702 4219 6704
rect 3620 6700 3626 6702
rect 4153 6699 4219 6702
rect 12157 6762 12223 6765
rect 12433 6762 12499 6765
rect 13629 6764 13695 6765
rect 13629 6762 13676 6764
rect 12157 6760 12499 6762
rect 12157 6704 12162 6760
rect 12218 6704 12438 6760
rect 12494 6704 12499 6760
rect 12157 6702 12499 6704
rect 13584 6760 13676 6762
rect 13584 6704 13634 6760
rect 13584 6702 13676 6704
rect 12157 6699 12223 6702
rect 12433 6699 12499 6702
rect 13629 6700 13676 6702
rect 13740 6700 13746 6764
rect 14181 6762 14247 6765
rect 17902 6762 17908 6764
rect 14181 6760 17908 6762
rect 14181 6704 14186 6760
rect 14242 6704 17908 6760
rect 14181 6702 17908 6704
rect 13629 6699 13695 6700
rect 14181 6699 14247 6702
rect 17902 6700 17908 6702
rect 17972 6700 17978 6764
rect 18413 6762 18479 6765
rect 19200 6762 20000 6792
rect 18413 6760 20000 6762
rect 18413 6704 18418 6760
rect 18474 6704 20000 6760
rect 18413 6702 20000 6704
rect 18413 6699 18479 6702
rect 19200 6672 20000 6702
rect 11697 6626 11763 6629
rect 12433 6626 12499 6629
rect 13721 6626 13787 6629
rect 11697 6624 13787 6626
rect 11697 6568 11702 6624
rect 11758 6568 12438 6624
rect 12494 6568 13726 6624
rect 13782 6568 13787 6624
rect 11697 6566 13787 6568
rect 11697 6563 11763 6566
rect 12433 6563 12499 6566
rect 13721 6563 13787 6566
rect 5394 6560 5710 6561
rect 0 6490 800 6520
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 14290 6495 14606 6496
rect 1853 6490 1919 6493
rect 0 6488 1919 6490
rect 0 6432 1858 6488
rect 1914 6432 1919 6488
rect 0 6430 1919 6432
rect 0 6400 800 6430
rect 1853 6427 1919 6430
rect 12249 6490 12315 6493
rect 12985 6490 13051 6493
rect 12249 6488 13051 6490
rect 12249 6432 12254 6488
rect 12310 6432 12990 6488
rect 13046 6432 13051 6488
rect 12249 6430 13051 6432
rect 12249 6427 12315 6430
rect 12985 6427 13051 6430
rect 4337 6354 4403 6357
rect 12157 6354 12223 6357
rect 4337 6352 12223 6354
rect 4337 6296 4342 6352
rect 4398 6296 12162 6352
rect 12218 6296 12223 6352
rect 4337 6294 12223 6296
rect 4337 6291 4403 6294
rect 12157 6291 12223 6294
rect 12801 6354 12867 6357
rect 14774 6354 14780 6356
rect 12801 6352 14780 6354
rect 12801 6296 12806 6352
rect 12862 6296 14780 6352
rect 12801 6294 14780 6296
rect 12801 6291 12867 6294
rect 14774 6292 14780 6294
rect 14844 6354 14850 6356
rect 18045 6354 18111 6357
rect 14844 6352 18111 6354
rect 14844 6296 18050 6352
rect 18106 6296 18111 6352
rect 14844 6294 18111 6296
rect 14844 6292 14850 6294
rect 18045 6291 18111 6294
rect 18413 6354 18479 6357
rect 19200 6354 20000 6384
rect 18413 6352 20000 6354
rect 18413 6296 18418 6352
rect 18474 6296 20000 6352
rect 18413 6294 20000 6296
rect 18413 6291 18479 6294
rect 19200 6264 20000 6294
rect 2221 6218 2287 6221
rect 5809 6218 5875 6221
rect 9070 6218 9076 6220
rect 2221 6216 9076 6218
rect 2221 6160 2226 6216
rect 2282 6160 5814 6216
rect 5870 6160 9076 6216
rect 2221 6158 9076 6160
rect 2221 6155 2287 6158
rect 5809 6155 5875 6158
rect 9070 6156 9076 6158
rect 9140 6156 9146 6220
rect 15653 6218 15719 6221
rect 18229 6218 18295 6221
rect 15653 6216 18295 6218
rect 15653 6160 15658 6216
rect 15714 6160 18234 6216
rect 18290 6160 18295 6216
rect 15653 6158 18295 6160
rect 15653 6155 15719 6158
rect 18229 6155 18295 6158
rect 0 6082 800 6112
rect 1485 6082 1551 6085
rect 0 6080 1551 6082
rect 0 6024 1490 6080
rect 1546 6024 1551 6080
rect 0 6022 1551 6024
rect 0 5992 800 6022
rect 1485 6019 1551 6022
rect 3601 6082 3667 6085
rect 4797 6082 4863 6085
rect 7373 6082 7439 6085
rect 3601 6080 7439 6082
rect 3601 6024 3606 6080
rect 3662 6024 4802 6080
rect 4858 6024 7378 6080
rect 7434 6024 7439 6080
rect 3601 6022 7439 6024
rect 3601 6019 3667 6022
rect 4797 6019 4863 6022
rect 7373 6019 7439 6022
rect 3170 6016 3486 6017
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 16514 5951 16830 5952
rect 4337 5946 4403 5949
rect 5165 5946 5231 5949
rect 4337 5944 5231 5946
rect 4337 5888 4342 5944
rect 4398 5888 5170 5944
rect 5226 5888 5231 5944
rect 4337 5886 5231 5888
rect 4337 5883 4403 5886
rect 5165 5883 5231 5886
rect 17033 5946 17099 5949
rect 19200 5946 20000 5976
rect 17033 5944 20000 5946
rect 17033 5888 17038 5944
rect 17094 5888 20000 5944
rect 17033 5886 20000 5888
rect 17033 5883 17099 5886
rect 19200 5856 20000 5886
rect 3141 5810 3207 5813
rect 3734 5810 3740 5812
rect 3141 5808 3740 5810
rect 3141 5752 3146 5808
rect 3202 5752 3740 5808
rect 3141 5750 3740 5752
rect 3141 5747 3207 5750
rect 3734 5748 3740 5750
rect 3804 5748 3810 5812
rect 4705 5810 4771 5813
rect 12249 5810 12315 5813
rect 16573 5810 16639 5813
rect 4705 5808 11898 5810
rect 4705 5752 4710 5808
rect 4766 5752 11898 5808
rect 4705 5750 11898 5752
rect 4705 5747 4771 5750
rect 0 5674 800 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 800 5614
rect 1577 5611 1643 5614
rect 3049 5674 3115 5677
rect 4153 5674 4219 5677
rect 3049 5672 4219 5674
rect 3049 5616 3054 5672
rect 3110 5616 4158 5672
rect 4214 5616 4219 5672
rect 3049 5614 4219 5616
rect 3049 5611 3115 5614
rect 4153 5611 4219 5614
rect 1669 5540 1735 5541
rect 1669 5536 1716 5540
rect 1780 5538 1786 5540
rect 3417 5538 3483 5541
rect 4708 5538 4768 5747
rect 6729 5674 6795 5677
rect 10593 5674 10659 5677
rect 11697 5674 11763 5677
rect 6729 5672 11763 5674
rect 6729 5616 6734 5672
rect 6790 5616 10598 5672
rect 10654 5616 11702 5672
rect 11758 5616 11763 5672
rect 6729 5614 11763 5616
rect 11838 5674 11898 5750
rect 12249 5808 16639 5810
rect 12249 5752 12254 5808
rect 12310 5752 16578 5808
rect 16634 5752 16639 5808
rect 12249 5750 16639 5752
rect 12249 5747 12315 5750
rect 16573 5747 16639 5750
rect 13302 5674 13308 5676
rect 11838 5614 13308 5674
rect 6729 5611 6795 5614
rect 10593 5611 10659 5614
rect 11697 5611 11763 5614
rect 13302 5612 13308 5614
rect 13372 5674 13378 5676
rect 13670 5674 13676 5676
rect 13372 5614 13676 5674
rect 13372 5612 13378 5614
rect 13670 5612 13676 5614
rect 13740 5612 13746 5676
rect 16021 5674 16087 5677
rect 17401 5674 17467 5677
rect 16021 5672 17467 5674
rect 16021 5616 16026 5672
rect 16082 5616 17406 5672
rect 17462 5616 17467 5672
rect 16021 5614 17467 5616
rect 16021 5611 16087 5614
rect 17401 5611 17467 5614
rect 1669 5480 1674 5536
rect 1669 5476 1716 5480
rect 1780 5478 1826 5538
rect 3417 5536 4768 5538
rect 3417 5480 3422 5536
rect 3478 5480 4768 5536
rect 3417 5478 4768 5480
rect 18413 5538 18479 5541
rect 19200 5538 20000 5568
rect 18413 5536 20000 5538
rect 18413 5480 18418 5536
rect 18474 5480 20000 5536
rect 18413 5478 20000 5480
rect 1780 5476 1786 5478
rect 1669 5475 1735 5476
rect 3417 5475 3483 5478
rect 18413 5475 18479 5478
rect 5394 5472 5710 5473
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 19200 5448 20000 5478
rect 14290 5407 14606 5408
rect 0 5266 800 5296
rect 1485 5266 1551 5269
rect 0 5264 1551 5266
rect 0 5208 1490 5264
rect 1546 5208 1551 5264
rect 0 5206 1551 5208
rect 0 5176 800 5206
rect 1485 5203 1551 5206
rect 2129 5266 2195 5269
rect 6729 5266 6795 5269
rect 2129 5264 6795 5266
rect 2129 5208 2134 5264
rect 2190 5208 6734 5264
rect 6790 5208 6795 5264
rect 2129 5206 6795 5208
rect 2129 5203 2195 5206
rect 6729 5203 6795 5206
rect 11145 5266 11211 5269
rect 17033 5268 17099 5269
rect 16982 5266 16988 5268
rect 11145 5264 16988 5266
rect 17052 5264 17099 5268
rect 11145 5208 11150 5264
rect 11206 5208 16988 5264
rect 17094 5208 17099 5264
rect 11145 5206 16988 5208
rect 11145 5203 11211 5206
rect 16982 5204 16988 5206
rect 17052 5204 17099 5208
rect 17033 5203 17099 5204
rect 4654 5068 4660 5132
rect 4724 5130 4730 5132
rect 7097 5130 7163 5133
rect 4724 5128 7163 5130
rect 4724 5072 7102 5128
rect 7158 5072 7163 5128
rect 4724 5070 7163 5072
rect 4724 5068 4730 5070
rect 7097 5067 7163 5070
rect 18505 5130 18571 5133
rect 19200 5130 20000 5160
rect 18505 5128 20000 5130
rect 18505 5072 18510 5128
rect 18566 5072 20000 5128
rect 18505 5070 20000 5072
rect 18505 5067 18571 5070
rect 19200 5040 20000 5070
rect 3170 4928 3486 4929
rect 0 4858 800 4888
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 16514 4863 16830 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 1945 4722 2011 4725
rect 6269 4722 6335 4725
rect 1945 4720 6746 4722
rect 1945 4664 1950 4720
rect 2006 4664 6274 4720
rect 6330 4664 6746 4720
rect 1945 4662 6746 4664
rect 1945 4659 2011 4662
rect 6269 4659 6335 4662
rect 6686 4586 6746 4662
rect 6862 4660 6868 4724
rect 6932 4722 6938 4724
rect 10133 4722 10199 4725
rect 6932 4720 10199 4722
rect 6932 4664 10138 4720
rect 10194 4664 10199 4720
rect 6932 4662 10199 4664
rect 6932 4660 6938 4662
rect 10133 4659 10199 4662
rect 16297 4722 16363 4725
rect 19200 4722 20000 4752
rect 16297 4720 20000 4722
rect 16297 4664 16302 4720
rect 16358 4664 20000 4720
rect 16297 4662 20000 4664
rect 16297 4659 16363 4662
rect 19200 4632 20000 4662
rect 10961 4586 11027 4589
rect 6686 4584 11027 4586
rect 6686 4528 10966 4584
rect 11022 4528 11027 4584
rect 6686 4526 11027 4528
rect 10961 4523 11027 4526
rect 0 4450 800 4480
rect 1485 4450 1551 4453
rect 0 4448 1551 4450
rect 0 4392 1490 4448
rect 1546 4392 1551 4448
rect 0 4390 1551 4392
rect 0 4360 800 4390
rect 1485 4387 1551 4390
rect 17585 4450 17651 4453
rect 17902 4450 17908 4452
rect 17585 4448 17908 4450
rect 17585 4392 17590 4448
rect 17646 4392 17908 4448
rect 17585 4390 17908 4392
rect 17585 4387 17651 4390
rect 17902 4388 17908 4390
rect 17972 4388 17978 4452
rect 5394 4384 5710 4385
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 14290 4319 14606 4320
rect 17033 4314 17099 4317
rect 19200 4314 20000 4344
rect 17033 4312 20000 4314
rect 17033 4256 17038 4312
rect 17094 4256 20000 4312
rect 17033 4254 20000 4256
rect 17033 4251 17099 4254
rect 19200 4224 20000 4254
rect 2630 4178 2636 4180
rect 2454 4118 2636 4178
rect 0 4042 800 4072
rect 1485 4042 1551 4045
rect 0 4040 1551 4042
rect 0 3984 1490 4040
rect 1546 3984 1551 4040
rect 0 3982 1551 3984
rect 0 3952 800 3982
rect 1485 3979 1551 3982
rect 1669 4042 1735 4045
rect 2454 4042 2514 4118
rect 2630 4116 2636 4118
rect 2700 4178 2706 4180
rect 6913 4178 6979 4181
rect 2700 4176 6979 4178
rect 2700 4120 6918 4176
rect 6974 4120 6979 4176
rect 2700 4118 6979 4120
rect 2700 4116 2706 4118
rect 6913 4115 6979 4118
rect 10593 4178 10659 4181
rect 10593 4176 16682 4178
rect 10593 4120 10598 4176
rect 10654 4120 16682 4176
rect 10593 4118 16682 4120
rect 10593 4115 10659 4118
rect 3049 4044 3115 4045
rect 1669 4040 2514 4042
rect 1669 3984 1674 4040
rect 1730 3984 2514 4040
rect 1669 3982 2514 3984
rect 1669 3979 1735 3982
rect 2998 3980 3004 4044
rect 3068 4042 3115 4044
rect 3068 4040 3160 4042
rect 3110 3984 3160 4040
rect 3068 3982 3160 3984
rect 3068 3980 3115 3982
rect 3918 3980 3924 4044
rect 3988 4042 3994 4044
rect 11145 4042 11211 4045
rect 3988 4040 11211 4042
rect 3988 3984 11150 4040
rect 11206 3984 11211 4040
rect 3988 3982 11211 3984
rect 3988 3980 3994 3982
rect 3049 3979 3115 3980
rect 11145 3979 11211 3982
rect 12341 4042 12407 4045
rect 14958 4042 14964 4044
rect 12341 4040 14964 4042
rect 12341 3984 12346 4040
rect 12402 3984 14964 4040
rect 12341 3982 14964 3984
rect 12341 3979 12407 3982
rect 14958 3980 14964 3982
rect 15028 3980 15034 4044
rect 16622 4042 16682 4118
rect 18597 4042 18663 4045
rect 16622 4040 18663 4042
rect 16622 3984 18602 4040
rect 18658 3984 18663 4040
rect 16622 3982 18663 3984
rect 18597 3979 18663 3982
rect 1894 3844 1900 3908
rect 1964 3906 1970 3908
rect 2037 3906 2103 3909
rect 1964 3904 2103 3906
rect 1964 3848 2042 3904
rect 2098 3848 2103 3904
rect 1964 3846 2103 3848
rect 1964 3844 1970 3846
rect 2037 3843 2103 3846
rect 13670 3844 13676 3908
rect 13740 3906 13746 3908
rect 16113 3906 16179 3909
rect 13740 3904 16179 3906
rect 13740 3848 16118 3904
rect 16174 3848 16179 3904
rect 13740 3846 16179 3848
rect 13740 3844 13746 3846
rect 16113 3843 16179 3846
rect 17217 3906 17283 3909
rect 19200 3906 20000 3936
rect 17217 3904 20000 3906
rect 17217 3848 17222 3904
rect 17278 3848 20000 3904
rect 17217 3846 20000 3848
rect 17217 3843 17283 3846
rect 3170 3840 3486 3841
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 19200 3816 20000 3846
rect 16514 3775 16830 3776
rect 0 3634 800 3664
rect 1853 3634 1919 3637
rect 0 3632 1919 3634
rect 0 3576 1858 3632
rect 1914 3576 1919 3632
rect 0 3574 1919 3576
rect 0 3544 800 3574
rect 1853 3571 1919 3574
rect 7414 3572 7420 3636
rect 7484 3634 7490 3636
rect 9397 3634 9463 3637
rect 7484 3632 9463 3634
rect 7484 3576 9402 3632
rect 9458 3576 9463 3632
rect 7484 3574 9463 3576
rect 7484 3572 7490 3574
rect 9397 3571 9463 3574
rect 17401 3634 17467 3637
rect 17718 3634 17724 3636
rect 17401 3632 17724 3634
rect 17401 3576 17406 3632
rect 17462 3576 17724 3632
rect 17401 3574 17724 3576
rect 17401 3571 17467 3574
rect 17718 3572 17724 3574
rect 17788 3572 17794 3636
rect 2589 3498 2655 3501
rect 11237 3498 11303 3501
rect 15377 3498 15443 3501
rect 2589 3496 15443 3498
rect 2589 3440 2594 3496
rect 2650 3440 11242 3496
rect 11298 3440 15382 3496
rect 15438 3440 15443 3496
rect 2589 3438 15443 3440
rect 2589 3435 2655 3438
rect 11237 3435 11303 3438
rect 15377 3435 15443 3438
rect 18413 3498 18479 3501
rect 19200 3498 20000 3528
rect 18413 3496 20000 3498
rect 18413 3440 18418 3496
rect 18474 3440 20000 3496
rect 18413 3438 20000 3440
rect 18413 3435 18479 3438
rect 19200 3408 20000 3438
rect 1117 3362 1183 3365
rect 4337 3362 4403 3365
rect 1117 3360 4403 3362
rect 1117 3304 1122 3360
rect 1178 3304 4342 3360
rect 4398 3304 4403 3360
rect 1117 3302 4403 3304
rect 1117 3299 1183 3302
rect 4337 3299 4403 3302
rect 5394 3296 5710 3297
rect 0 3226 800 3256
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 14290 3231 14606 3232
rect 1485 3226 1551 3229
rect 0 3224 1551 3226
rect 0 3168 1490 3224
rect 1546 3168 1551 3224
rect 0 3166 1551 3168
rect 0 3136 800 3166
rect 1485 3163 1551 3166
rect 3417 3090 3483 3093
rect 4102 3090 4108 3092
rect 3417 3088 4108 3090
rect 3417 3032 3422 3088
rect 3478 3032 4108 3088
rect 3417 3030 4108 3032
rect 3417 3027 3483 3030
rect 4102 3028 4108 3030
rect 4172 3028 4178 3092
rect 6085 3090 6151 3093
rect 13997 3090 14063 3093
rect 6085 3088 14063 3090
rect 6085 3032 6090 3088
rect 6146 3032 14002 3088
rect 14058 3032 14063 3088
rect 6085 3030 14063 3032
rect 6085 3027 6151 3030
rect 13997 3027 14063 3030
rect 18045 3090 18111 3093
rect 19200 3090 20000 3120
rect 18045 3088 20000 3090
rect 18045 3032 18050 3088
rect 18106 3032 20000 3088
rect 18045 3030 20000 3032
rect 18045 3027 18111 3030
rect 19200 3000 20000 3030
rect 4337 2954 4403 2957
rect 8109 2954 8175 2957
rect 12617 2954 12683 2957
rect 4337 2952 12683 2954
rect 4337 2896 4342 2952
rect 4398 2896 8114 2952
rect 8170 2896 12622 2952
rect 12678 2896 12683 2952
rect 4337 2894 12683 2896
rect 4337 2891 4403 2894
rect 0 2818 800 2848
rect 4846 2821 4906 2894
rect 8109 2891 8175 2894
rect 12617 2891 12683 2894
rect 1577 2818 1643 2821
rect 0 2816 1643 2818
rect 0 2760 1582 2816
rect 1638 2760 1643 2816
rect 0 2758 1643 2760
rect 0 2728 800 2758
rect 1577 2755 1643 2758
rect 2037 2818 2103 2821
rect 2037 2816 2882 2818
rect 2037 2760 2042 2816
rect 2098 2760 2882 2816
rect 2037 2758 2882 2760
rect 2037 2755 2103 2758
rect 2822 2546 2882 2758
rect 4797 2816 4906 2821
rect 4797 2760 4802 2816
rect 4858 2760 4906 2816
rect 4797 2758 4906 2760
rect 4797 2755 4863 2758
rect 3170 2752 3486 2753
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 16514 2687 16830 2688
rect 3877 2684 3943 2685
rect 3877 2682 3924 2684
rect 3558 2680 3924 2682
rect 3988 2682 3994 2684
rect 13721 2682 13787 2685
rect 17493 2684 17559 2685
rect 14038 2682 14044 2684
rect 3558 2624 3882 2680
rect 3558 2622 3924 2624
rect 3558 2546 3618 2622
rect 3877 2620 3924 2622
rect 3988 2622 4034 2682
rect 13721 2680 14044 2682
rect 13721 2624 13726 2680
rect 13782 2624 14044 2680
rect 13721 2622 14044 2624
rect 3988 2620 3994 2622
rect 3877 2619 3943 2620
rect 13721 2619 13787 2622
rect 14038 2620 14044 2622
rect 14108 2620 14114 2684
rect 17493 2680 17540 2684
rect 17604 2682 17610 2684
rect 17769 2682 17835 2685
rect 19200 2682 20000 2712
rect 17493 2624 17498 2680
rect 17493 2620 17540 2624
rect 17604 2622 17650 2682
rect 17769 2680 20000 2682
rect 17769 2624 17774 2680
rect 17830 2624 20000 2680
rect 17769 2622 20000 2624
rect 17604 2620 17610 2622
rect 17493 2619 17559 2620
rect 17769 2619 17835 2622
rect 19200 2592 20000 2622
rect 2822 2486 3618 2546
rect 8150 2484 8156 2548
rect 8220 2546 8226 2548
rect 9397 2546 9463 2549
rect 8220 2544 9463 2546
rect 8220 2488 9402 2544
rect 9458 2488 9463 2544
rect 8220 2486 9463 2488
rect 8220 2484 8226 2486
rect 9397 2483 9463 2486
rect 0 2410 800 2440
rect 1853 2410 1919 2413
rect 0 2408 1919 2410
rect 0 2352 1858 2408
rect 1914 2352 1919 2408
rect 0 2350 1919 2352
rect 0 2320 800 2350
rect 1853 2347 1919 2350
rect 16941 2274 17007 2277
rect 19200 2274 20000 2304
rect 16941 2272 20000 2274
rect 16941 2216 16946 2272
rect 17002 2216 20000 2272
rect 16941 2214 20000 2216
rect 16941 2211 17007 2214
rect 5394 2208 5710 2209
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 19200 2184 20000 2214
rect 14290 2143 14606 2144
rect 0 2002 800 2032
rect 2221 2002 2287 2005
rect 0 2000 2287 2002
rect 0 1944 2226 2000
rect 2282 1944 2287 2000
rect 0 1942 2287 1944
rect 0 1912 800 1942
rect 2221 1939 2287 1942
rect 15837 1866 15903 1869
rect 19200 1866 20000 1896
rect 15837 1864 20000 1866
rect 15837 1808 15842 1864
rect 15898 1808 20000 1864
rect 15837 1806 20000 1808
rect 15837 1803 15903 1806
rect 19200 1776 20000 1806
rect 0 1594 800 1624
rect 2681 1594 2747 1597
rect 0 1592 2747 1594
rect 0 1536 2686 1592
rect 2742 1536 2747 1592
rect 0 1534 2747 1536
rect 0 1504 800 1534
rect 2681 1531 2747 1534
rect 15377 1458 15443 1461
rect 19200 1458 20000 1488
rect 15377 1456 20000 1458
rect 15377 1400 15382 1456
rect 15438 1400 20000 1456
rect 15377 1398 20000 1400
rect 15377 1395 15443 1398
rect 19200 1368 20000 1398
rect 0 1186 800 1216
rect 1945 1186 2011 1189
rect 0 1184 2011 1186
rect 0 1128 1950 1184
rect 2006 1128 2011 1184
rect 0 1126 2011 1128
rect 0 1096 800 1126
rect 1945 1123 2011 1126
rect 15193 1050 15259 1053
rect 19200 1050 20000 1080
rect 15193 1048 20000 1050
rect 15193 992 15198 1048
rect 15254 992 20000 1048
rect 15193 990 20000 992
rect 15193 987 15259 990
rect 19200 960 20000 990
rect 0 778 800 808
rect 1669 778 1735 781
rect 0 776 1735 778
rect 0 720 1674 776
rect 1730 720 1735 776
rect 0 718 1735 720
rect 0 688 800 718
rect 1669 715 1735 718
rect 15929 642 15995 645
rect 19200 642 20000 672
rect 15929 640 20000 642
rect 15929 584 15934 640
rect 15990 584 20000 640
rect 15929 582 20000 584
rect 15929 579 15995 582
rect 19200 552 20000 582
rect 0 370 800 400
rect 3785 370 3851 373
rect 0 368 3851 370
rect 0 312 3790 368
rect 3846 312 3851 368
rect 0 310 3851 312
rect 0 280 800 310
rect 3785 307 3851 310
<< via3 >>
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 3556 13908 3620 13972
rect 13492 13832 13556 13836
rect 13492 13776 13542 13832
rect 13542 13776 13556 13832
rect 13492 13772 13556 13776
rect 13676 13772 13740 13836
rect 17540 13772 17604 13836
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 3740 13560 3804 13564
rect 3740 13504 3790 13560
rect 3790 13504 3804 13560
rect 3740 13500 3804 13504
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 3924 12820 3988 12884
rect 6316 12880 6380 12884
rect 6316 12824 6366 12880
rect 6366 12824 6380 12880
rect 6316 12820 6380 12824
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 1716 12412 1780 12476
rect 14964 12412 15028 12476
rect 13860 12276 13924 12340
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 13492 11868 13556 11932
rect 9076 11460 9140 11524
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 5028 11324 5092 11388
rect 5212 11052 5276 11116
rect 7420 11052 7484 11116
rect 9260 11112 9324 11116
rect 9260 11056 9274 11112
rect 9274 11056 9324 11112
rect 9260 11052 9324 11056
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3924 10840 3988 10844
rect 3924 10784 3974 10840
rect 3974 10784 3988 10840
rect 3924 10780 3988 10784
rect 2820 10644 2884 10708
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 6500 10372 6564 10436
rect 16988 10372 17052 10436
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 5948 10236 6012 10300
rect 16068 10236 16132 10300
rect 4476 9964 4540 10028
rect 16068 10024 16132 10028
rect 16068 9968 16118 10024
rect 16118 9968 16132 10024
rect 16068 9964 16132 9968
rect 16988 9888 17052 9892
rect 16988 9832 17038 9888
rect 17038 9832 17052 9888
rect 16988 9828 17052 9832
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 3004 9692 3068 9756
rect 4108 9692 4172 9756
rect 6868 9692 6932 9756
rect 8156 9692 8220 9756
rect 14044 9752 14108 9756
rect 14044 9696 14058 9752
rect 14058 9696 14108 9752
rect 14044 9692 14108 9696
rect 17908 9752 17972 9756
rect 17908 9696 17922 9752
rect 17922 9696 17972 9752
rect 17908 9692 17972 9696
rect 3740 9420 3804 9484
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 4660 9420 4724 9484
rect 5948 9420 6012 9484
rect 13492 9284 13556 9348
rect 14780 9344 14844 9348
rect 14780 9288 14830 9344
rect 14830 9288 14844 9344
rect 14780 9284 14844 9288
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 4476 9012 4540 9076
rect 2452 8936 2516 8940
rect 2452 8880 2466 8936
rect 2466 8880 2516 8936
rect 2452 8876 2516 8880
rect 1900 8740 1964 8804
rect 5028 8740 5092 8804
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 13860 8604 13924 8668
rect 6500 8256 6564 8260
rect 6500 8200 6550 8256
rect 6550 8200 6564 8256
rect 6500 8196 6564 8200
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 5212 7516 5276 7580
rect 3740 7380 3804 7444
rect 6316 7380 6380 7444
rect 9260 7380 9324 7444
rect 2452 7244 2516 7308
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 17724 7032 17788 7036
rect 17724 6976 17774 7032
rect 17774 6976 17788 7032
rect 17724 6972 17788 6976
rect 3556 6700 3620 6764
rect 13676 6760 13740 6764
rect 13676 6704 13690 6760
rect 13690 6704 13740 6760
rect 13676 6700 13740 6704
rect 17908 6700 17972 6764
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 14780 6292 14844 6356
rect 9076 6156 9140 6220
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 3740 5748 3804 5812
rect 1716 5536 1780 5540
rect 13308 5612 13372 5676
rect 13676 5612 13740 5676
rect 1716 5480 1730 5536
rect 1730 5480 1780 5536
rect 1716 5476 1780 5480
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 16988 5264 17052 5268
rect 16988 5208 17038 5264
rect 17038 5208 17052 5264
rect 16988 5204 17052 5208
rect 4660 5068 4724 5132
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 6868 4660 6932 4724
rect 17908 4388 17972 4452
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 2636 4116 2700 4180
rect 3004 4040 3068 4044
rect 3004 3984 3054 4040
rect 3054 3984 3068 4040
rect 3004 3980 3068 3984
rect 3924 3980 3988 4044
rect 14964 3980 15028 4044
rect 1900 3844 1964 3908
rect 13676 3844 13740 3908
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 7420 3572 7484 3636
rect 17724 3572 17788 3636
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 4108 3028 4172 3092
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 3924 2680 3988 2684
rect 3924 2624 3938 2680
rect 3938 2624 3988 2680
rect 3924 2620 3988 2624
rect 14044 2620 14108 2684
rect 17540 2680 17604 2684
rect 17540 2624 17554 2680
rect 17554 2624 17604 2680
rect 17540 2620 17604 2624
rect 8156 2484 8220 2548
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 3555 13972 3621 13973
rect 3555 13908 3556 13972
rect 3620 13908 3621 13972
rect 3555 13907 3621 13908
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 1715 12476 1781 12477
rect 1715 12412 1716 12476
rect 1780 12412 1781 12476
rect 1715 12411 1781 12412
rect 1718 5541 1778 12411
rect 3168 11456 3488 12480
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 2819 10708 2885 10709
rect 2819 10644 2820 10708
rect 2884 10644 2885 10708
rect 2819 10643 2885 10644
rect 2451 8940 2517 8941
rect 2451 8876 2452 8940
rect 2516 8876 2517 8940
rect 2451 8875 2517 8876
rect 1899 8804 1965 8805
rect 1899 8740 1900 8804
rect 1964 8740 1965 8804
rect 1899 8739 1965 8740
rect 1715 5540 1781 5541
rect 1715 5476 1716 5540
rect 1780 5476 1781 5540
rect 1715 5475 1781 5476
rect 1902 3909 1962 8739
rect 2454 7309 2514 8875
rect 2451 7308 2517 7309
rect 2451 7244 2452 7308
rect 2516 7244 2517 7308
rect 2451 7243 2517 7244
rect 2822 6930 2882 10643
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3003 9756 3069 9757
rect 3003 9692 3004 9756
rect 3068 9692 3069 9756
rect 3003 9691 3069 9692
rect 2638 6870 2882 6930
rect 2638 4181 2698 6870
rect 2635 4180 2701 4181
rect 2635 4116 2636 4180
rect 2700 4116 2701 4180
rect 2635 4115 2701 4116
rect 3006 4045 3066 9691
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 6016 3488 7040
rect 3558 6765 3618 13907
rect 3739 13564 3805 13565
rect 3739 13500 3740 13564
rect 3804 13500 3805 13564
rect 3739 13499 3805 13500
rect 3742 9485 3802 13499
rect 5392 13088 5712 14112
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 3926 10845 3986 12819
rect 5392 12000 5712 13024
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 6315 12884 6381 12885
rect 6315 12820 6316 12884
rect 6380 12820 6381 12884
rect 6315 12819 6381 12820
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5027 11388 5093 11389
rect 5027 11324 5028 11388
rect 5092 11324 5093 11388
rect 5027 11323 5093 11324
rect 3923 10844 3989 10845
rect 3923 10780 3924 10844
rect 3988 10780 3989 10844
rect 3923 10779 3989 10780
rect 4475 10028 4541 10029
rect 4475 9964 4476 10028
rect 4540 9964 4541 10028
rect 4475 9963 4541 9964
rect 4107 9756 4173 9757
rect 4107 9692 4108 9756
rect 4172 9692 4173 9756
rect 4107 9691 4173 9692
rect 3739 9484 3805 9485
rect 3739 9420 3740 9484
rect 3804 9420 3805 9484
rect 3739 9419 3805 9420
rect 3739 7444 3805 7445
rect 3739 7380 3740 7444
rect 3804 7380 3805 7444
rect 3739 7379 3805 7380
rect 3555 6764 3621 6765
rect 3555 6700 3556 6764
rect 3620 6700 3621 6764
rect 3555 6699 3621 6700
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 4928 3488 5952
rect 3742 5813 3802 7379
rect 3739 5812 3805 5813
rect 3739 5748 3740 5812
rect 3804 5748 3805 5812
rect 3739 5747 3805 5748
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3003 4044 3069 4045
rect 3003 3980 3004 4044
rect 3068 3980 3069 4044
rect 3003 3979 3069 3980
rect 1899 3908 1965 3909
rect 1899 3844 1900 3908
rect 1964 3844 1965 3908
rect 1899 3843 1965 3844
rect 3168 3840 3488 4864
rect 3923 4044 3989 4045
rect 3923 3980 3924 4044
rect 3988 3980 3989 4044
rect 3923 3979 3989 3980
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 3926 2685 3986 3979
rect 4110 3093 4170 9691
rect 4478 9077 4538 9963
rect 4659 9484 4725 9485
rect 4659 9420 4660 9484
rect 4724 9420 4725 9484
rect 4659 9419 4725 9420
rect 4475 9076 4541 9077
rect 4475 9012 4476 9076
rect 4540 9012 4541 9076
rect 4475 9011 4541 9012
rect 4662 5133 4722 9419
rect 5030 8805 5090 11323
rect 5211 11116 5277 11117
rect 5211 11052 5212 11116
rect 5276 11052 5277 11116
rect 5211 11051 5277 11052
rect 5027 8804 5093 8805
rect 5027 8740 5028 8804
rect 5092 8740 5093 8804
rect 5027 8739 5093 8740
rect 5214 7581 5274 11051
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5947 10300 6013 10301
rect 5947 10236 5948 10300
rect 6012 10236 6013 10300
rect 5947 10235 6013 10236
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 5950 9485 6010 10235
rect 5947 9484 6013 9485
rect 5947 9420 5948 9484
rect 6012 9420 6013 9484
rect 5947 9419 6013 9420
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5211 7580 5277 7581
rect 5211 7516 5212 7580
rect 5276 7516 5277 7580
rect 5211 7515 5277 7516
rect 5392 6560 5712 7584
rect 6318 7445 6378 12819
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 11456 7936 12480
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9075 11524 9141 11525
rect 9075 11460 9076 11524
rect 9140 11460 9141 11524
rect 9075 11459 9141 11460
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 6499 10436 6565 10437
rect 6499 10372 6500 10436
rect 6564 10372 6565 10436
rect 6499 10371 6565 10372
rect 6502 8261 6562 10371
rect 6867 9756 6933 9757
rect 6867 9692 6868 9756
rect 6932 9692 6933 9756
rect 6867 9691 6933 9692
rect 6499 8260 6565 8261
rect 6499 8196 6500 8260
rect 6564 8196 6565 8260
rect 6499 8195 6565 8196
rect 6315 7444 6381 7445
rect 6315 7380 6316 7444
rect 6380 7380 6381 7444
rect 6315 7379 6381 7380
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 4659 5132 4725 5133
rect 4659 5068 4660 5132
rect 4724 5068 4725 5132
rect 4659 5067 4725 5068
rect 5392 4384 5712 5408
rect 6870 4725 6930 9691
rect 6867 4724 6933 4725
rect 6867 4660 6868 4724
rect 6932 4660 6933 4724
rect 6867 4659 6933 4660
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 7422 3637 7482 11051
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7419 3636 7485 3637
rect 7419 3572 7420 3636
rect 7484 3572 7485 3636
rect 7419 3571 7485 3572
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 4107 3092 4173 3093
rect 4107 3028 4108 3092
rect 4172 3028 4173 3092
rect 4107 3027 4173 3028
rect 3923 2684 3989 2685
rect 3923 2620 3924 2684
rect 3988 2620 3989 2684
rect 3923 2619 3989 2620
rect 5392 2208 5712 3232
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2752 7936 3776
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2128 7936 2688
rect 8158 2549 8218 9691
rect 9078 6221 9138 11459
rect 9259 11116 9325 11117
rect 9259 11052 9260 11116
rect 9324 11052 9325 11116
rect 9259 11051 9325 11052
rect 9262 7445 9322 11051
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9259 7444 9325 7445
rect 9259 7380 9260 7444
rect 9324 7380 9325 7444
rect 9259 7379 9325 7380
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9075 6220 9141 6221
rect 9075 6156 9076 6220
rect 9140 6156 9141 6220
rect 9075 6155 9141 6156
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 8155 2548 8221 2549
rect 8155 2484 8156 2548
rect 8220 2484 8221 2548
rect 8155 2483 8221 2484
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 13491 13836 13557 13837
rect 13491 13772 13492 13836
rect 13556 13772 13557 13836
rect 13491 13771 13557 13772
rect 13675 13836 13741 13837
rect 13675 13772 13676 13836
rect 13740 13772 13741 13836
rect 13675 13771 13741 13772
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 13494 12450 13554 13771
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 13310 12390 13554 12450
rect 13310 5677 13370 12390
rect 13491 11932 13557 11933
rect 13491 11868 13492 11932
rect 13556 11868 13557 11932
rect 13491 11867 13557 11868
rect 13494 9349 13554 11867
rect 13491 9348 13557 9349
rect 13491 9284 13492 9348
rect 13556 9284 13557 9348
rect 13491 9283 13557 9284
rect 13678 6765 13738 13771
rect 14288 13088 14608 14112
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 13859 12340 13925 12341
rect 13859 12276 13860 12340
rect 13924 12276 13925 12340
rect 13859 12275 13925 12276
rect 13862 8669 13922 12275
rect 14288 12000 14608 13024
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16512 13632 16832 14656
rect 17539 13836 17605 13837
rect 17539 13772 17540 13836
rect 17604 13772 17605 13836
rect 17539 13771 17605 13772
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 14963 12476 15029 12477
rect 14963 12412 14964 12476
rect 15028 12412 15029 12476
rect 14963 12411 15029 12412
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14043 9756 14109 9757
rect 14043 9692 14044 9756
rect 14108 9692 14109 9756
rect 14043 9691 14109 9692
rect 13859 8668 13925 8669
rect 13859 8604 13860 8668
rect 13924 8604 13925 8668
rect 13859 8603 13925 8604
rect 13675 6764 13741 6765
rect 13675 6700 13676 6764
rect 13740 6700 13741 6764
rect 13675 6699 13741 6700
rect 13307 5676 13373 5677
rect 13307 5612 13308 5676
rect 13372 5612 13373 5676
rect 13307 5611 13373 5612
rect 13675 5676 13741 5677
rect 13675 5612 13676 5676
rect 13740 5612 13741 5676
rect 13675 5611 13741 5612
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 13678 3909 13738 5611
rect 13675 3908 13741 3909
rect 13675 3844 13676 3908
rect 13740 3844 13741 3908
rect 13675 3843 13741 3844
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14046 2685 14106 9691
rect 14288 8736 14608 9760
rect 14779 9348 14845 9349
rect 14779 9284 14780 9348
rect 14844 9284 14845 9348
rect 14779 9283 14845 9284
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14782 6357 14842 9283
rect 14779 6356 14845 6357
rect 14779 6292 14780 6356
rect 14844 6292 14845 6356
rect 14779 6291 14845 6292
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 14966 4045 15026 12411
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16987 10436 17053 10437
rect 16987 10372 16988 10436
rect 17052 10372 17053 10436
rect 16987 10371 17053 10372
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16067 10300 16133 10301
rect 16067 10236 16068 10300
rect 16132 10236 16133 10300
rect 16067 10235 16133 10236
rect 16070 10029 16130 10235
rect 16067 10028 16133 10029
rect 16067 9964 16068 10028
rect 16132 9964 16133 10028
rect 16067 9963 16133 9964
rect 16512 9280 16832 10304
rect 16990 9893 17050 10371
rect 16987 9892 17053 9893
rect 16987 9828 16988 9892
rect 17052 9828 17053 9892
rect 16987 9827 17053 9828
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16990 5269 17050 9827
rect 16987 5268 17053 5269
rect 16987 5204 16988 5268
rect 17052 5204 17053 5268
rect 16987 5203 17053 5204
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 14963 4044 15029 4045
rect 14963 3980 14964 4044
rect 15028 3980 15029 4044
rect 14963 3979 15029 3980
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14043 2684 14109 2685
rect 14043 2620 14044 2684
rect 14108 2620 14109 2684
rect 14043 2619 14109 2620
rect 14288 2208 14608 3232
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 3840 16832 4864
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
rect 17542 2685 17602 13771
rect 17907 9756 17973 9757
rect 17907 9692 17908 9756
rect 17972 9692 17973 9756
rect 17907 9691 17973 9692
rect 17723 7036 17789 7037
rect 17723 6972 17724 7036
rect 17788 6972 17789 7036
rect 17723 6971 17789 6972
rect 17726 3637 17786 6971
rect 17910 6765 17970 9691
rect 17907 6764 17973 6765
rect 17907 6700 17908 6764
rect 17972 6700 17973 6764
rect 17907 6699 17973 6700
rect 17910 4453 17970 6699
rect 17907 4452 17973 4453
rect 17907 4388 17908 4452
rect 17972 4388 17973 4452
rect 17907 4387 17973 4388
rect 17723 3636 17789 3637
rect 17723 3572 17724 3636
rect 17788 3572 17789 3636
rect 17723 3571 17789 3572
rect 17539 2684 17605 2685
rect 17539 2620 17540 2684
rect 17604 2620 17605 2684
rect 17539 2619 17605 2620
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform -1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 2760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 2300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform -1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform -1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 17112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform 1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform -1 0 16560 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 6532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 7084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3864 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5152 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 2852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 13984 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 15364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 14996 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 16560 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 11960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 18584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6440 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1649977179
transform -1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 1932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 5980 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform -1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater114_A
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1649977179
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1649977179
transform 1 0 10488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_131
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_17
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_59
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_87
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_75
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_51
timestamp 1649977179
transform 1 0 5796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1649977179
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_86
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_58
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_96
timestamp 1649977179
transform 1 0 9936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_122
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_95
timestamp 1649977179
transform 1 0 9844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_168
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_95
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_16
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_47
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_116
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1649977179
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_31
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_53
timestamp 1649977179
transform 1 0 5980 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_122
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_178
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_113
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_152
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_170
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_32
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_96
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_141
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp 1649977179
transform 1 0 15548 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_55
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_79
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_91
timestamp 1649977179
transform 1 0 9476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1649977179
transform 1 0 6164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_76
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_101
timestamp 1649977179
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _34_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform 1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 12144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 17848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 4968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform -1 0 3220 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform -1 0 3588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 3220 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1649977179
transform -1 0 4692 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform -1 0 2300 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1649977179
transform -1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 17296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1649977179
transform -1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 16560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1649977179
transform -1 0 18584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15272 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10488 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 15088 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13432 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7912 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8096 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10580 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7544 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5796 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9844 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8188 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7268 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6532 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8096 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13524 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12880 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11592 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14904 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15180 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_ipin_0.mux_l2_in_3__132 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3864 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5336 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_0.mux_l2_in_3__133
timestamp 1649977179
transform -1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2760 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_1.mux_l2_in_3__134
timestamp 1649977179
transform -1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_2.mux_l2_in_3__141
timestamp 1649977179
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_3.mux_l2_in_3__142
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3128 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3496 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7268 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_4.mux_l2_in_3__126
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5520 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4692 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_5.mux_l2_in_3__127
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4784 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_6.mux_l2_in_3__128
timestamp 1649977179
transform -1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5980 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_7.mux_l2_in_3__129
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6256 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7268 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_8.mux_l2_in_3__130
timestamp 1649977179
transform -1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_9.mux_l2_in_3__131
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_10.mux_l2_in_3__135
timestamp 1649977179
transform 1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform -1 0 16468 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5612 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_11.mux_l2_in_3__136
timestamp 1649977179
transform -1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15364 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_12.mux_l2_in_3__137
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_13.mux_l2_in_3__138
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_14.mux_l2_in_3__139
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18032 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17112 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_15.mux_l2_in_3__140
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16376 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output47 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 16284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 10396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 17296 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 12144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 16744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output108
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater110
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater111
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater112
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater113
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater114
timestamp 1649977179
transform -1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater115
timestamp 1649977179
transform -1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater116
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater117
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater118
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater119
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater120
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater121
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater122
timestamp 1649977179
transform 1 0 10488 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater123
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater124
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater125
timestamp 1649977179
transform -1 0 3680 0 -1 11968
box -38 -48 314 592
<< labels >>
flabel metal2 s 1122 16400 1178 17200 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 1 nsew signal input
flabel metal2 s 3330 16400 3386 17200 0 FreeSans 224 90 0 0 SC_IN_TOP
port 2 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 3 nsew signal tristate
flabel metal2 s 5538 16400 5594 17200 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 4 nsew signal tristate
flabel metal4 s 5392 2128 5712 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 7616 2128 7936 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 12064 2128 12384 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 16512 2128 16832 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 bottom_grid_pin_0_
port 7 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 bottom_grid_pin_10_
port 8 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 bottom_grid_pin_11_
port 9 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 bottom_grid_pin_12_
port 10 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 bottom_grid_pin_13_
port 11 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 bottom_grid_pin_14_
port 12 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 bottom_grid_pin_15_
port 13 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 bottom_grid_pin_1_
port 14 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_grid_pin_2_
port 15 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 bottom_grid_pin_3_
port 16 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 bottom_grid_pin_4_
port 17 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 bottom_grid_pin_5_
port 18 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 bottom_grid_pin_6_
port 19 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 bottom_grid_pin_7_
port 20 nsew signal tristate
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 bottom_grid_pin_8_
port 21 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 bottom_grid_pin_9_
port 22 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_0_
port 23 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_1_lower
port 24 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_1_upper
port 25 nsew signal tristate
flabel metal2 s 7746 16400 7802 17200 0 FreeSans 224 90 0 0 ccff_head
port 26 nsew signal input
flabel metal2 s 9954 16400 10010 17200 0 FreeSans 224 90 0 0 ccff_tail
port 27 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 28 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 29 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 30 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 31 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 32 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 33 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 34 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 35 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 36 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 37 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 38 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 39 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 40 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 41 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 42 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 43 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 44 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 45 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 46 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 47 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 48 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 49 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 50 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 51 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 52 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 53 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 54 nsew signal tristate
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 55 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 56 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 57 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 58 nsew signal tristate
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 59 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 60 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 61 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 62 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 63 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 64 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 65 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 66 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 67 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 68 nsew signal input
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 69 nsew signal input
flabel metal3 s 19200 13200 20000 13320 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 70 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 71 nsew signal input
flabel metal3 s 19200 14016 20000 14136 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 72 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 73 nsew signal input
flabel metal3 s 19200 14832 20000 14952 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 74 nsew signal input
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 75 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 76 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 77 nsew signal input
flabel metal3 s 19200 16464 20000 16584 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 78 nsew signal input
flabel metal3 s 19200 9120 20000 9240 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 79 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 80 nsew signal input
flabel metal3 s 19200 9936 20000 10056 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 81 nsew signal input
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 82 nsew signal input
flabel metal3 s 19200 10752 20000 10872 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 83 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 84 nsew signal input
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 85 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 86 nsew signal input
flabel metal3 s 19200 12384 20000 12504 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 87 nsew signal input
flabel metal3 s 19200 552 20000 672 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 88 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 89 nsew signal tristate
flabel metal3 s 19200 5040 20000 5160 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 90 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 91 nsew signal tristate
flabel metal3 s 19200 5856 20000 5976 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 92 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 93 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 94 nsew signal tristate
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 95 nsew signal tristate
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 96 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 97 nsew signal tristate
flabel metal3 s 19200 8304 20000 8424 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 98 nsew signal tristate
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 99 nsew signal tristate
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 100 nsew signal tristate
flabel metal3 s 19200 1776 20000 1896 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 101 nsew signal tristate
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 102 nsew signal tristate
flabel metal3 s 19200 2592 20000 2712 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 103 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 104 nsew signal tristate
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 105 nsew signal tristate
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 106 nsew signal tristate
flabel metal3 s 19200 4224 20000 4344 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 107 nsew signal tristate
flabel metal2 s 14370 16400 14426 17200 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 108 nsew signal tristate
flabel metal2 s 16578 16400 16634 17200 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 109 nsew signal input
flabel metal2 s 18786 16400 18842 17200 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 110 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 111 nsew signal input
flabel metal3 s 0 280 800 400 0 FreeSans 480 0 0 0 prog_clk_0_W_out
port 112 nsew signal tristate
flabel metal2 s 12162 16400 12218 17200 0 FreeSans 224 90 0 0 top_grid_pin_0_
port 113 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
